/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
main
**
**
**
*****************************************************************************/
module
main(
InstDone,
Jen,
Jin,
Jout,
R1,
R10,
R11,
R12,
R13,
R14,
R15,
R16,
R17,
R18,
R19,
R2,
R20,
R21,
R22,
R23,
R24,
R25,
R26,
R27,
R28,
R29,
R3,
R30,
R31,
R4,
R5,
R6,
R7,
R8,
R9,
clk,
nop,
rst
);
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
Jen;
input
[31:0]
Jin;
input
clk;
input
rst;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
InstDone;
output
[31:0]
Jout;
output
[31:0]
R1;
output
[31:0]
R10;
output
[31:0]
R11;
output
[31:0]
R12;
output
[31:0]
R13;
output
[31:0]
R14;
output
[31:0]
R15;
output
[31:0]
R16;
output
[31:0]
R17;
output
[31:0]
R18;
output
[31:0]
R19;
output
[31:0]
R2;
output
[31:0]
R20;
output
[31:0]
R21;
output
[31:0]
R22;
output
[31:0]
R23;
output
[31:0]
R24;
output
[31:0]
R25;
output
[31:0]
R26;
output
[31:0]
R27;
output
[31:0]
R28;
output
[31:0]
R29;
output
[31:0]
R3;
output
[31:0]
R30;
output
[31:0]
R31;
output
[31:0]
R4;
output
[31:0]
R5;
output
[31:0]
R6;
output
[31:0]
R7;
output
[31:0]
R8;
output
[31:0]
R9;
output
nop;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
[31:0]
s_logisimBus0;
wire
[4:0]
s_logisimBus10;
wire
[31:0]
s_logisimBus13;
wire
[15:0]
s_logisimBus14;
wire
[4:0]
s_logisimBus15;
wire
[31:0]
s_logisimBus16;
wire
[8:0]
s_logisimBus17;
wire
[31:0]
s_logisimBus18;
wire
[5:0]
s_logisimBus19;
wire
[31:0]
s_logisimBus22;
wire
[31:0]
s_logisimBus23;
wire
[4:0]
s_logisimBus24;
wire
[31:0]
s_logisimBus25;
wire
[8:0]
s_logisimBus26;
wire
[4:0]
s_logisimBus27;
wire
[31:0]
s_logisimBus28;
wire
[31:0]
s_logisimBus29;
wire
[8:0]
s_logisimBus3;
wire
[8:0]
s_logisimBus30;
wire
[31:0]
s_logisimBus32;
wire
[31:0]
s_logisimBus35;
wire
[31:0]
s_logisimBus36;
wire
[31:0]
s_logisimBus37;
wire
[4:0]
s_logisimBus38;
wire
[8:0]
s_logisimBus39;
wire
[3:0]
s_logisimBus4;
wire
[31:0]
s_logisimBus45;
wire
[4:0]
s_logisimBus46;
wire
[8:0]
s_logisimBus47;
wire
[5:0]
s_logisimBus5;
wire
[31:0]
s_logisimBus50;
wire
[31:0]
s_logisimBus54;
wire
[31:0]
s_logisimBus55;
wire
[31:0]
s_logisimBus56;
wire
[31:0]
s_logisimBus57;
wire
[31:0]
s_logisimBus58;
wire
[31:0]
s_logisimBus59;
wire
[4:0]
s_logisimBus6;
wire
[31:0]
s_logisimBus60;
wire
[31:0]
s_logisimBus61;
wire
[31:0]
s_logisimBus62;
wire
[31:0]
s_logisimBus63;
wire
[31:0]
s_logisimBus64;
wire
[31:0]
s_logisimBus65;
wire
[31:0]
s_logisimBus66;
wire
[31:0]
s_logisimBus67;
wire
[31:0]
s_logisimBus68;
wire
[31:0]
s_logisimBus69;
wire
[31:0]
s_logisimBus70;
wire
[31:0]
s_logisimBus71;
wire
[31:0]
s_logisimBus72;
wire
[31:0]
s_logisimBus73;
wire
[31:0]
s_logisimBus74;
wire
[31:0]
s_logisimBus75;
wire
[31:0]
s_logisimBus76;
wire
[31:0]
s_logisimBus77;
wire
[31:0]
s_logisimBus78;
wire
[31:0]
s_logisimBus79;
wire
[31:0]
s_logisimBus8;
wire
[31:0]
s_logisimBus80;
wire
[31:0]
s_logisimBus81;
wire
[31:0]
s_logisimBus82;
wire
[31:0]
s_logisimBus83;
wire
[31:0]
s_logisimBus84;
wire
[31:0]
s_logisimBus85;
wire
[31:0]
s_logisimBus86;
wire
s_logisimNet1;
wire
s_logisimNet11;
wire
s_logisimNet12;
wire
s_logisimNet2;
wire
s_logisimNet20;
wire
s_logisimNet21;
wire
s_logisimNet33;
wire
s_logisimNet34;
wire
s_logisimNet40;
wire
s_logisimNet41;
wire
s_logisimNet42;
wire
s_logisimNet43;
wire
s_logisimNet44;
wire
s_logisimNet48;
wire
s_logisimNet51;
wire
s_logisimNet52;
wire
s_logisimNet53;
wire
s_logisimNet7;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
all
input
connections
are
defined
**
*******************************************************************************/
assign
s_logisimBus45[31:0]
=
Jin;
assign
s_logisimNet12
=
rst;
assign
s_logisimNet2
=
Jen;
assign
s_logisimNet43
=
clk;
/*******************************************************************************
**
Here
all
output
connections
are
defined
**
*******************************************************************************/
assign
InstDone
=
s_logisimNet11;
assign
Jout
=
s_logisimBus29[31:0];
assign
R1
=
s_logisimBus56[31:0];
assign
R10
=
s_logisimBus65[31:0];
assign
R11
=
s_logisimBus66[31:0];
assign
R12
=
s_logisimBus67[31:0];
assign
R13
=
s_logisimBus68[31:0];
assign
R14
=
s_logisimBus69[31:0];
assign
R15
=
s_logisimBus70[31:0];
assign
R16
=
s_logisimBus71[31:0];
assign
R17
=
s_logisimBus72[31:0];
assign
R18
=
s_logisimBus73[31:0];
assign
R19
=
s_logisimBus74[31:0];
assign
R2
=
s_logisimBus57[31:0];
assign
R20
=
s_logisimBus75[31:0];
assign
R21
=
s_logisimBus76[31:0];
assign
R22
=
s_logisimBus77[31:0];
assign
R23
=
s_logisimBus78[31:0];
assign
R24
=
s_logisimBus79[31:0];
assign
R25
=
s_logisimBus80[31:0];
assign
R26
=
s_logisimBus81[31:0];
assign
R27
=
s_logisimBus82[31:0];
assign
R28
=
s_logisimBus83[31:0];
assign
R29
=
s_logisimBus84[31:0];
assign
R3
=
s_logisimBus58[31:0];
assign
R30
=
s_logisimBus85[31:0];
assign
R31
=
s_logisimBus86[31:0];
assign
R4
=
s_logisimBus59[31:0];
assign
R5
=
s_logisimBus60[31:0];
assign
R6
=
s_logisimBus61[31:0];
assign
R7
=
s_logisimBus62[31:0];
assign
R8
=
s_logisimBus63[31:0];
assign
R9
=
s_logisimBus64[31:0];
assign
nop
=
s_logisimNet41;
/*******************************************************************************
**
Here
all
in-lined
components
are
defined
**
*******************************************************************************/
assign
s_logisimBus13[0]
=
s_logisimBus10[0];
assign
s_logisimBus13[1]
=
s_logisimBus10[1];
assign
s_logisimBus13[2]
=
s_logisimBus10[2];
assign
s_logisimBus13[3]
=
s_logisimBus10[3];
assign
s_logisimBus13[4]
=
s_logisimBus10[4];
assign
s_logisimBus13[5]
=
1'b0;
assign
s_logisimBus13[6]
=
1'b0;
assign
s_logisimBus13[7]
=
1'b0;
assign
s_logisimBus13[8]
=
1'b0;
assign
s_logisimBus13[9]
=
1'b0;
assign
s_logisimBus13[10]
=
1'b0;
assign
s_logisimBus13[11]
=
1'b0;
assign
s_logisimBus13[12]
=
1'b0;
assign
s_logisimBus13[13]
=
1'b0;
assign
s_logisimBus13[14]
=
1'b0;
assign
s_logisimBus13[15]
=
1'b0;
assign
s_logisimBus13[16]
=
1'b0;
assign
s_logisimBus13[17]
=
1'b0;
assign
s_logisimBus13[18]
=
1'b0;
assign
s_logisimBus13[19]
=
1'b0;
assign
s_logisimBus13[20]
=
1'b0;
assign
s_logisimBus13[21]
=
1'b0;
assign
s_logisimBus13[22]
=
1'b0;
assign
s_logisimBus13[23]
=
1'b0;
assign
s_logisimBus13[24]
=
1'b0;
assign
s_logisimBus13[25]
=
1'b0;
assign
s_logisimBus13[26]
=
1'b0;
assign
s_logisimBus13[27]
=
1'b0;
assign
s_logisimBus13[28]
=
1'b0;
assign
s_logisimBus13[29]
=
1'b0;
assign
s_logisimBus13[30]
=
1'b0;
assign
s_logisimBus13[31]
=
1'b0;
assign
s_logisimBus47[8:0]
=
{1'b0,
8'h01};
assign
s_logisimBus46[4:0]
=
{1'b0,
4'h0};
assign
s_logisimBus32[0]
=
s_logisimBus14[0];
assign
s_logisimBus32[1]
=
s_logisimBus14[1];
assign
s_logisimBus32[2]
=
s_logisimBus14[2];
assign
s_logisimBus32[3]
=
s_logisimBus14[3];
assign
s_logisimBus32[4]
=
s_logisimBus14[4];
assign
s_logisimBus32[5]
=
s_logisimBus14[5];
assign
s_logisimBus32[6]
=
s_logisimBus14[6];
assign
s_logisimBus32[7]
=
s_logisimBus14[7];
assign
s_logisimBus32[8]
=
s_logisimBus14[8];
assign
s_logisimBus32[9]
=
s_logisimBus14[9];
assign
s_logisimBus32[10]
=
s_logisimBus14[10];
assign
s_logisimBus32[11]
=
s_logisimBus14[11];
assign
s_logisimBus32[12]
=
s_logisimBus14[12];
assign
s_logisimBus32[13]
=
s_logisimBus14[13];
assign
s_logisimBus32[14]
=
s_logisimBus14[14];
assign
s_logisimBus32[15]
=
s_logisimBus14[15];
assign
s_logisimBus32[16]
=
s_logisimBus14[15];
assign
s_logisimBus32[17]
=
s_logisimBus14[15];
assign
s_logisimBus32[18]
=
s_logisimBus14[15];
assign
s_logisimBus32[19]
=
s_logisimBus14[15];
assign
s_logisimBus32[20]
=
s_logisimBus14[15];
assign
s_logisimBus32[21]
=
s_logisimBus14[15];
assign
s_logisimBus32[22]
=
s_logisimBus14[15];
assign
s_logisimBus32[23]
=
s_logisimBus14[15];
assign
s_logisimBus32[24]
=
s_logisimBus14[15];
assign
s_logisimBus32[25]
=
s_logisimBus14[15];
assign
s_logisimBus32[26]
=
s_logisimBus14[15];
assign
s_logisimBus32[27]
=
s_logisimBus14[15];
assign
s_logisimBus32[28]
=
s_logisimBus14[15];
assign
s_logisimBus32[29]
=
s_logisimBus14[15];
assign
s_logisimBus32[30]
=
s_logisimBus14[15];
assign
s_logisimBus32[31]
=
s_logisimBus14[15];
/*******************************************************************************
**
Here
all
normal
components
are
defined
**
*******************************************************************************/
AND_GATE
#(.BubblesMask(2'b01))
GATES_1
(.input1(s_logisimNet33),
.input2(s_logisimNet52),
.result(s_logisimNet40));
AND_GATE
#(.BubblesMask(2'b10))
GATES_2
(.input1(s_logisimNet43),
.input2(s_logisimNet41),
.result(s_logisimNet48));
Multiplexer_bus_2
#(.nrOfBits(32))
PLEXERS_3
(.enable(1'b1),
.muxIn_0(s_logisimBus18[31:0]),
.muxIn_1(s_logisimBus13[31:0]),
.muxOut(s_logisimBus37[31:0]),
.sel(s_logisimNet7));
Multiplexer_bus_2
#(.nrOfBits(32))
PLEXERS_4
(.enable(1'b1),
.muxIn_0(s_logisimBus54[31:0]),
.muxIn_1(s_logisimBus55[31:0]),
.muxOut(s_logisimBus8[31:0]),
.sel(s_logisimNet7));
Multiplexer_bus_2
#(.nrOfBits(9))
PLEXERS_5
(.enable(1'b1),
.muxIn_0(s_logisimBus3[8:0]),
.muxIn_1(s_logisimBus39[8:0]),
.muxOut(s_logisimBus30[8:0]),
.sel(s_logisimNet40));
Multiplexer_bus_2
#(.nrOfBits(9))
PLEXERS_6
(.enable(1'b1),
.muxIn_0(s_logisimBus30[8:0]),
.muxIn_1(s_logisimBus14[8:0]),
.muxOut(s_logisimBus26[8:0]),
.sel(s_logisimNet44));
Multiplexer_bus_2
#(.nrOfBits(5))
PLEXERS_7
(.enable(1'b1),
.muxIn_0(s_logisimBus27[4:0]),
.muxIn_1(s_logisimBus38[4:0]),
.muxOut(s_logisimBus15[4:0]),
.sel(s_logisimNet42));
Multiplexer_bus_2
#(.nrOfBits(32))
PLEXERS_8
(.enable(1'b1),
.muxIn_0(s_logisimBus36[31:0]),
.muxIn_1(s_logisimBus50[31:0]),
.muxOut(s_logisimBus0[31:0]),
.sel(s_logisimNet34));
Multiplexer_bus_2
#(.nrOfBits(32))
PLEXERS_9
(.enable(1'b1),
.muxIn_0(s_logisimBus0[31:0]),
.muxIn_1(s_logisimBus35[31:0]),
.muxOut(s_logisimBus16[31:0]),
.sel(s_logisimNet21));
Multiplexer_bus_2
#(.nrOfBits(5))
PLEXERS_10
(.enable(1'b1),
.muxIn_0(s_logisimBus46[4:0]),
.muxIn_1(s_logisimBus15[4:0]),
.muxOut(s_logisimBus6[4:0]),
.sel(s_logisimNet20));
Multiplexer_bus_2
#(.nrOfBits(32))
PLEXERS_11
(.enable(1'b1),
.muxIn_0(s_logisimBus55[31:0]),
.muxIn_1(s_logisimBus32[31:0]),
.muxOut(s_logisimBus18[31:0]),
.sel(s_logisimNet1));
Adder
#(.extendedBits(10),
.nrOfBits(9))
ARITH_12
(.carryIn(1'b0),
.carryOut(),
.dataA(s_logisimBus3[8:0]),
.dataB(s_logisimBus32[8:0]),
.result(s_logisimBus39[8:0]));
Adder
#(.extendedBits(10),
.nrOfBits(9))
ARITH_13
(.carryIn(1'b0),
.carryOut(),
.dataA(s_logisimBus17[8:0]),
.dataB(s_logisimBus47[8:0]),
.result(s_logisimBus3[8:0]));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(9))
pc
(.clock(s_logisimNet48),
.clockEnable(1'b1),
.d(s_logisimBus26[8:0]),
.q(s_logisimBus17[8:0]),
.reset(s_logisimNet12),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(32))
HI
(.clock(s_logisimNet48),
.clockEnable(s_logisimNet53),
.d(s_logisimBus25[31:0]),
.q(s_logisimBus35[31:0]),
.reset(1'b0),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(32))
LO
(.clock(s_logisimNet48),
.clockEnable(s_logisimNet53),
.d(s_logisimBus36[31:0]),
.q(s_logisimBus23[31:0]),
.reset(1'b0),
.tick(1'b1));
/*******************************************************************************
**
Here
all
sub-circuits
are
defined
**
*******************************************************************************/
jtag_ram512
Dmem
(.Addr(s_logisimBus36[8:0]),
.Din(s_logisimBus55[31:0]),
.Dout(s_logisimBus50[31:0]),
.Jen(s_logisimNet2),
.Jin(s_logisimBus22[31:0]),
.Jout(s_logisimBus29[31:0]),
.Wen(s_logisimNet51),
.clk(s_logisimNet48));
ALU
x3
(.InstDone(s_logisimNet11),
.a(s_logisimBus8[31:0]),
.aluop(s_logisimBus4[3:0]),
.b(s_logisimBus37[31:0]),
.clk(s_logisimNet43),
.res_high(s_logisimBus25[31:0]),
.res_low(s_logisimBus36[31:0]),
.zero(s_logisimNet33));
InstructionDecode
x1
(.Instruction(s_logisimBus28[31:0]),
.func(s_logisimBus19[5:0]),
.imm(s_logisimBus14[15:0]),
.opCode(s_logisimBus5[5:0]),
.rd(s_logisimBus38[4:0]),
.rs(s_logisimBus27[4:0]),
.rt(s_logisimBus24[4:0]),
.shmt(s_logisimBus10[4:0]));
ControlUnit
ControlUnit_1
(.ALUop(s_logisimBus4[3:0]),
.ALUsrc(s_logisimNet1),
.Rtype(),
.branch(s_logisimNet52),
.divv(s_logisimNet53),
.func(s_logisimBus19[5:0]),
.inst(s_logisimNet11),
.j(s_logisimNet44),
.main_clock(s_logisimNet43),
.memRead(),
.memToReg(s_logisimNet34),
.memWrite(s_logisimNet51),
.mohi(s_logisimNet21),
.nop(s_logisimNet41),
.opCode(s_logisimBus5[5:0]),
.regDst(s_logisimNet42),
.regWrite(s_logisimNet20),
.shmt(s_logisimNet7));
jtag_ram512
Imem
(.Addr(s_logisimBus17[8:0]),
.Din(32'd0),
.Dout(s_logisimBus28[31:0]),
.Jen(s_logisimNet2),
.Jin(s_logisimBus45[31:0]),
.Jout(s_logisimBus22[31:0]),
.Wen(1'b0),
.clk(s_logisimNet48));
regfile
x4
(.Aread0(s_logisimBus24[4:0]),
.Aread1(s_logisimBus27[4:0]),
.Awrite(s_logisimBus6[4:0]),
.Dread0(s_logisimBus54[31:0]),
.Dread1(s_logisimBus55[31:0]),
.Dwrite(s_logisimBus16[31:0]),
.R1(s_logisimBus56[31:0]),
.R10(s_logisimBus65[31:0]),
.R11(s_logisimBus66[31:0]),
.R12(s_logisimBus67[31:0]),
.R13(s_logisimBus68[31:0]),
.R14(s_logisimBus69[31:0]),
.R15(s_logisimBus70[31:0]),
.R16(s_logisimBus71[31:0]),
.R17(s_logisimBus72[31:0]),
.R18(s_logisimBus73[31:0]),
.R19(s_logisimBus74[31:0]),
.R2(s_logisimBus57[31:0]),
.R20(s_logisimBus75[31:0]),
.R21(s_logisimBus76[31:0]),
.R22(s_logisimBus77[31:0]),
.R23(s_logisimBus78[31:0]),
.R24(s_logisimBus79[31:0]),
.R25(s_logisimBus80[31:0]),
.R26(s_logisimBus81[31:0]),
.R27(s_logisimBus82[31:0]),
.R28(s_logisimBus83[31:0]),
.R29(s_logisimBus84[31:0]),
.R3(s_logisimBus58[31:0]),
.R30(s_logisimBus85[31:0]),
.R31(s_logisimBus86[31:0]),
.R4(s_logisimBus59[31:0]),
.R5(s_logisimBus60[31:0]),
.R6(s_logisimBus61[31:0]),
.R7(s_logisimBus62[31:0]),
.R8(s_logisimBus63[31:0]),
.R9(s_logisimBus64[31:0]),
.clk(s_logisimNet48),
.rst(s_logisimNet12));
endmodule