/******************************************************************************
 ** Logisim-evolution goes FPGA automatic generated Verilog code             **
 ** https://github.com/logisim-evolution/                                    **
 **                                                                          **
 ** Component : SLTI                                                         **
 **                                                                          **
 *****************************************************************************/

module SLTI( a,
             b,
             res_low );

   /*******************************************************************************
   ** The inputs are defined here                                                **
   *******************************************************************************/
   input [31:0] a;
   input [31:0] b;

   /*******************************************************************************
   ** The outputs are defined here                                               **
   *******************************************************************************/
   output [31:0] res_low;

   /*******************************************************************************
   ** The wires are defined here                                                 **
   *******************************************************************************/
   wire [31:0] s_logisimBus1;
   wire [31:0] s_logisimBus2;
   wire [31:0] s_logisimBus3;
   wire        s_logisimNet0;

   /*******************************************************************************
   ** The module functionality is described here                                 **
   *******************************************************************************/

   /*******************************************************************************
   ** Here all input connections are defined                                     **
   *******************************************************************************/
   assign s_logisimBus2[31:0] = a;
   assign s_logisimBus3[31:0] = b;

   /*******************************************************************************
   ** Here all output connections are defined                                    **
   *******************************************************************************/
   assign res_low = s_logisimBus1[31:0];

   /*******************************************************************************
   ** Here all in-lined components are defined                                   **
   *******************************************************************************/

   // Bit Extender
   assign  s_logisimBus1[0]  =  s_logisimNet0;
   assign  s_logisimBus1[1]  =  1'b0;
   assign  s_logisimBus1[2]  =  1'b0;
   assign  s_logisimBus1[3]  =  1'b0;
   assign  s_logisimBus1[4]  =  1'b0;
   assign  s_logisimBus1[5]  =  1'b0;
   assign  s_logisimBus1[6]  =  1'b0;
   assign  s_logisimBus1[7]  =  1'b0;
   assign  s_logisimBus1[8]  =  1'b0;
   assign  s_logisimBus1[9]  =  1'b0;
   assign  s_logisimBus1[10]  =  1'b0;
   assign  s_logisimBus1[11]  =  1'b0;
   assign  s_logisimBus1[12]  =  1'b0;
   assign  s_logisimBus1[13]  =  1'b0;
   assign  s_logisimBus1[14]  =  1'b0;
   assign  s_logisimBus1[15]  =  1'b0;
   assign  s_logisimBus1[16]  =  1'b0;
   assign  s_logisimBus1[17]  =  1'b0;
   assign  s_logisimBus1[18]  =  1'b0;
   assign  s_logisimBus1[19]  =  1'b0;
   assign  s_logisimBus1[20]  =  1'b0;
   assign  s_logisimBus1[21]  =  1'b0;
   assign  s_logisimBus1[22]  =  1'b0;
   assign  s_logisimBus1[23]  =  1'b0;
   assign  s_logisimBus1[24]  =  1'b0;
   assign  s_logisimBus1[25]  =  1'b0;
   assign  s_logisimBus1[26]  =  1'b0;
   assign  s_logisimBus1[27]  =  1'b0;
   assign  s_logisimBus1[28]  =  1'b0;
   assign  s_logisimBus1[29]  =  1'b0;
   assign  s_logisimBus1[30]  =  1'b0;
   assign  s_logisimBus1[31]  =  1'b0;


   /*******************************************************************************
   ** Here all normal components are defined                                     **
   *******************************************************************************/
   Comparator #(.nrOfBits(32),
                .twosComplement(1))
      ARITH_1 (.aEqualsB(),
               .aGreaterThanB(),
               .aLessThanB(s_logisimNet0),
               .dataA(s_logisimBus2[31:0]),
               .dataB(s_logisimBus3[31:0]));


endmodule
