/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
SRAA
**
**
**
*****************************************************************************/
module
SRAA(
a,
b,
res_high,
res_low
);
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
[31:0]
a;
input
[31:0]
b;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
[31:0]
res_high;
output
[31:0]
res_low;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
[31:0]
s_logisimBus0;
wire
[31:0]
s_logisimBus1;
wire
[31:0]
s_logisimBus10;
wire
[31:0]
s_logisimBus11;
wire
[31:0]
s_logisimBus2;
wire
[31:0]
s_logisimBus3;
wire
[31:0]
s_logisimBus4;
wire
[31:0]
s_logisimBus5;
wire
[31:0]
s_logisimBus6;
wire
[31:0]
s_logisimBus8;
wire
[31:0]
s_logisimBus9;
wire
s_logisimNet12;
wire
s_logisimNet7;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
all
input
connections
are
defined
**
*******************************************************************************/
assign
s_logisimBus0[31:0]
=
b;
assign
s_logisimBus2[31:0]
=
a;
/*******************************************************************************
**
Here
all
output
connections
are
defined
**
*******************************************************************************/
assign
res_high
=
s_logisimBus11[31:0];
assign
res_low
=
s_logisimBus1[31:0];
/*******************************************************************************
**
Here
all
in-lined
components
are
defined
**
*******************************************************************************/
assign
s_logisimBus9[0]
=
s_logisimBus2[31];
assign
s_logisimBus9[1]
=
s_logisimBus2[31];
assign
s_logisimBus9[2]
=
s_logisimBus2[31];
assign
s_logisimBus9[3]
=
s_logisimBus2[31];
assign
s_logisimBus9[4]
=
s_logisimBus2[31];
assign
s_logisimBus9[5]
=
s_logisimBus2[31];
assign
s_logisimBus9[6]
=
s_logisimBus2[31];
assign
s_logisimBus9[7]
=
s_logisimBus2[31];
assign
s_logisimBus9[8]
=
s_logisimBus2[31];
assign
s_logisimBus9[9]
=
s_logisimBus2[31];
assign
s_logisimBus9[10]
=
s_logisimBus2[31];
assign
s_logisimBus9[11]
=
s_logisimBus2[31];
assign
s_logisimBus9[12]
=
s_logisimBus2[31];
assign
s_logisimBus9[13]
=
s_logisimBus2[31];
assign
s_logisimBus9[14]
=
s_logisimBus2[31];
assign
s_logisimBus9[15]
=
s_logisimBus2[31];
assign
s_logisimBus9[16]
=
s_logisimBus2[31];
assign
s_logisimBus9[17]
=
s_logisimBus2[31];
assign
s_logisimBus9[18]
=
s_logisimBus2[31];
assign
s_logisimBus9[19]
=
s_logisimBus2[31];
assign
s_logisimBus9[20]
=
s_logisimBus2[31];
assign
s_logisimBus9[21]
=
s_logisimBus2[31];
assign
s_logisimBus9[22]
=
s_logisimBus2[31];
assign
s_logisimBus9[23]
=
s_logisimBus2[31];
assign
s_logisimBus9[24]
=
s_logisimBus2[31];
assign
s_logisimBus9[25]
=
s_logisimBus2[31];
assign
s_logisimBus9[26]
=
s_logisimBus2[31];
assign
s_logisimBus9[27]
=
s_logisimBus2[31];
assign
s_logisimBus9[28]
=
s_logisimBus2[31];
assign
s_logisimBus9[29]
=
s_logisimBus2[31];
assign
s_logisimBus9[30]
=
s_logisimBus2[31];
assign
s_logisimBus9[31]
=
s_logisimBus2[31];
assign
s_logisimBus10[31:0]
=
32'h00000020;
assign
s_logisimBus5[31:0]
=
32'h0000001F;
assign
s_logisimBus11[0]
=
s_logisimBus1[31];
assign
s_logisimBus11[1]
=
s_logisimBus1[31];
assign
s_logisimBus11[2]
=
s_logisimBus1[31];
assign
s_logisimBus11[3]
=
s_logisimBus1[31];
assign
s_logisimBus11[4]
=
s_logisimBus1[31];
assign
s_logisimBus11[5]
=
s_logisimBus1[31];
assign
s_logisimBus11[6]
=
s_logisimBus1[31];
assign
s_logisimBus11[7]
=
s_logisimBus1[31];
assign
s_logisimBus11[8]
=
s_logisimBus1[31];
assign
s_logisimBus11[9]
=
s_logisimBus1[31];
assign
s_logisimBus11[10]
=
s_logisimBus1[31];
assign
s_logisimBus11[11]
=
s_logisimBus1[31];
assign
s_logisimBus11[12]
=
s_logisimBus1[31];
assign
s_logisimBus11[13]
=
s_logisimBus1[31];
assign
s_logisimBus11[14]
=
s_logisimBus1[31];
assign
s_logisimBus11[15]
=
s_logisimBus1[31];
assign
s_logisimBus11[16]
=
s_logisimBus1[31];
assign
s_logisimBus11[17]
=
s_logisimBus1[31];
assign
s_logisimBus11[18]
=
s_logisimBus1[31];
assign
s_logisimBus11[19]
=
s_logisimBus1[31];
assign
s_logisimBus11[20]
=
s_logisimBus1[31];
assign
s_logisimBus11[21]
=
s_logisimBus1[31];
assign
s_logisimBus11[22]
=
s_logisimBus1[31];
assign
s_logisimBus11[23]
=
s_logisimBus1[31];
assign
s_logisimBus11[24]
=
s_logisimBus1[31];
assign
s_logisimBus11[25]
=
s_logisimBus1[31];
assign
s_logisimBus11[26]
=
s_logisimBus1[31];
assign
s_logisimBus11[27]
=
s_logisimBus1[31];
assign
s_logisimBus11[28]
=
s_logisimBus1[31];
assign
s_logisimBus11[29]
=
s_logisimBus1[31];
assign
s_logisimBus11[30]
=
s_logisimBus1[31];
assign
s_logisimBus11[31]
=
s_logisimBus1[31];
/*******************************************************************************
**
Here
all
normal
components
are
defined
**
*******************************************************************************/
AND_GATE_BUS
#(.BubblesMask(2'b00),
.NrOfBits(32))
GATES_1
(.input1(s_logisimBus0[31:0]),
.input2(s_logisimBus5[31:0]),
.result(s_logisimBus8[31:0]));
OR_GATE_BUS
#(.BubblesMask(2'b00),
.NrOfBits(32))
GATES_2
(.input1(s_logisimBus3[31:0]),
.input2(s_logisimBus4[31:0]),
.result(s_logisimBus1[31:0]));
Subtractor
#(.extendedBits(33),
.nrOfBits(32))
ARITH_3
(.borrowIn(1'b0),
.borrowOut(),
.dataA(s_logisimBus10[31:0]),
.dataB(s_logisimBus8[31:0]),
.result(s_logisimBus6[31:0]));
/*******************************************************************************
**
Here
all
sub-circuits
are
defined
**
*******************************************************************************/
SRLL
sth1
(.a(s_logisimBus2[31:0]),
.b(s_logisimBus0[31:0]),
.res_high(),
.res_low(s_logisimBus3[31:0]));
SLLL
sth2
(.a(s_logisimBus9[31:0]),
.b(s_logisimBus6[31:0]),
.res_high(),
.res_low(s_logisimBus4[31:0]));
endmodule