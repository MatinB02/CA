/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
InstructionDecode
**
**
**
*****************************************************************************/
module
InstructionDecode(
Instruction,
func,
imm,
opCode,
rd,
rs,
rt,
shmt
);
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
[31:0]
Instruction;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
[5:0]
func;
output
[15:0]
imm;
output
[5:0]
opCode;
output
[4:0]
rd;
output
[4:0]
rs;
output
[4:0]
rt;
output
[4:0]
shmt;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
[31:0]
s_logisimBus1;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
all
input
connections
are
defined
**
*******************************************************************************/
assign
s_logisimBus1[31:0]
=
Instruction;
/*******************************************************************************
**
Here
all
output
connections
are
defined
**
*******************************************************************************/
assign
func
=
s_logisimBus1[5:0];
assign
imm
=
s_logisimBus1[15:0];
assign
opCode
=
s_logisimBus1[31:26];
assign
rd
=
s_logisimBus1[15:11];
assign
rs
=
s_logisimBus1[20:16];
assign
rt
=
s_logisimBus1[25:21];
assign
shmt
=
s_logisimBus1[10:6];
endmodule