/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
main
**
**
**
*****************************************************************************/
module
main(
clk,
in1,
load,
out1
);
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
clk;
input
[31:0]
in1;
input
load;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
[31:0]
out1;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
[31:0]
s_logisimBus0;
wire
[31:0]
s_logisimBus2;
wire
[31:0]
s_logisimBus3;
wire
[31:0]
s_logisimBus4;
wire
[31:0]
s_logisimBus5;
wire
[31:0]
s_logisimBus6;
wire
[31:0]
s_logisimBus7;
wire
s_logisimNet1;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
all
input
connections
are
defined
**
*******************************************************************************/
assign
s_logisimBus4[31:0]
=
in1;
assign
s_logisimNet1
=
clk;
/*******************************************************************************
**
Here
all
output
connections
are
defined
**
*******************************************************************************/
assign
out1
=
s_logisimBus7[31:0];
/*******************************************************************************
**
Here
all
normal
components
are
defined
**
*******************************************************************************/
AND_GATE_BUS
#(.BubblesMask(2'b00),
.NrOfBits(32))
GATES_1
(.input1(s_logisimBus3[31:0]),
.input2(s_logisimBus4[31:0]),
.result(s_logisimBus5[31:0]));
Negator
#(.nrOfBits(32))
ARITH_2
(.dataX(s_logisimBus4[31:0]),
.minDataX(s_logisimBus0[31:0]));
Negator
#(.nrOfBits(32))
ARITH_3
(.dataX(s_logisimBus2[31:0]),
.minDataX(s_logisimBus6[31:0]));
Adder
#(.extendedBits(33),
.nrOfBits(32))
ARITH_4
(.carryIn(1'b0),
.carryOut(),
.dataA(s_logisimBus6[31:0]),
.dataB(s_logisimBus4[31:0]),
.result(s_logisimBus7[31:0]));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(32))
MEMORY_5
(.clock(s_logisimNet1),
.clockEnable(1'b1),
.d(s_logisimBus0[31:0]),
.q(s_logisimBus3[31:0]),
.reset(1'b0),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(32))
MEMORY_6
(.clock(s_logisimNet1),
.clockEnable(1'b1),
.d(s_logisimBus5[31:0]),
.q(s_logisimBus2[31:0]),
.reset(1'b0),
.tick(1'b1));
endmodule