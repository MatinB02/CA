/******************************************************************************
 ** Logisim-evolution goes FPGA automatic generated Verilog code             **
 ** https://github.com/logisim-evolution/                                    **
 **                                                                          **
 ** Component : SRL_fadd                                                     **
 **                                                                          **
 *****************************************************************************/

module SRL_fadd( a,
                 b,
                 one_signal,
                 res_low );

   /*******************************************************************************
   ** The inputs are defined here                                                **
   *******************************************************************************/
   input [31:0] a;
   input [31:0] b;

   /*******************************************************************************
   ** The outputs are defined here                                               **
   *******************************************************************************/
   output        one_signal;
   output [31:0] res_low;

   /*******************************************************************************
   ** The wires are defined here                                                 **
   *******************************************************************************/
   wire [31:0] s_logisimBus0;
   wire [31:0] s_logisimBus1;
   wire [31:0] s_logisimBus10;
   wire [31:0] s_logisimBus12;
   wire [31:0] s_logisimBus13;
   wire [31:0] s_logisimBus16;
   wire [31:0] s_logisimBus19;
   wire [31:0] s_logisimBus20;
   wire [4:0]  s_logisimBus22;
   wire [31:0] s_logisimBus29;
   wire [31:0] s_logisimBus3;
   wire [4:0]  s_logisimBus30;
   wire [4:0]  s_logisimBus31;
   wire [31:0] s_logisimBus4;
   wire [31:0] s_logisimBus8;
   wire [31:0] s_logisimBus9;
   wire        s_logisimNet11;
   wire        s_logisimNet14;
   wire        s_logisimNet15;
   wire        s_logisimNet17;
   wire        s_logisimNet18;
   wire        s_logisimNet2;
   wire        s_logisimNet21;
   wire        s_logisimNet23;
   wire        s_logisimNet24;
   wire        s_logisimNet25;
   wire        s_logisimNet26;
   wire        s_logisimNet27;
   wire        s_logisimNet28;
   wire        s_logisimNet5;
   wire        s_logisimNet6;
   wire        s_logisimNet7;

   /*******************************************************************************
   ** The module functionality is described here                                 **
   *******************************************************************************/

   /*******************************************************************************
   ** Here all wiring is defined                                                 **
   *******************************************************************************/
   assign s_logisimBus22[0] = s_logisimNet24;
   assign s_logisimBus22[1] = s_logisimNet25;
   assign s_logisimBus22[2] = s_logisimNet26;
   assign s_logisimBus22[3] = s_logisimNet27;
   assign s_logisimBus22[4] = s_logisimNet28;
   assign s_logisimBus30[0] = s_logisimNet6;
   assign s_logisimBus30[1] = s_logisimNet5;
   assign s_logisimBus30[2] = s_logisimNet2;
   assign s_logisimBus30[3] = s_logisimNet11;
   assign s_logisimBus30[4] = s_logisimNet18;
   assign s_logisimNet11    = s_logisimBus9[3];
   assign s_logisimNet18    = s_logisimBus9[4];
   assign s_logisimNet2     = s_logisimBus9[2];
   assign s_logisimNet24    = s_logisimBus4[0];
   assign s_logisimNet25    = s_logisimBus4[1];
   assign s_logisimNet26    = s_logisimBus4[2];
   assign s_logisimNet27    = s_logisimBus4[3];
   assign s_logisimNet28    = s_logisimBus4[4];
   assign s_logisimNet5     = s_logisimBus9[1];
   assign s_logisimNet6     = s_logisimBus9[0];

   /*******************************************************************************
   ** Here all input connections are defined                                     **
   *******************************************************************************/
   assign s_logisimBus0[31:0] = a;
   assign s_logisimBus9[31:0] = b;

   /*******************************************************************************
   ** Here all output connections are defined                                    **
   *******************************************************************************/
   assign one_signal = s_logisimNet15;
   assign res_low    = s_logisimBus3[31:0];

   /*******************************************************************************
   ** Here all in-lined components are defined                                   **
   *******************************************************************************/

   // Constant
   assign  s_logisimBus29[31:0]  =  32'h00000001;


   // Constant
   assign  s_logisimBus10[31:0]  =  32'h00000000;


   // Constant
   assign  s_logisimBus1[31:0]  =  32'h0000001F;


   // Constant
   assign  s_logisimBus31[4:0]  =  {1'b0, 4'h1};


   // Constant
   assign  s_logisimBus20[31:0]  =  32'h00000000;


   // NOT Gate
   assign s_logisimNet14 = ~s_logisimNet7;

   /*******************************************************************************
   ** Here all normal components are defined                                     **
   *******************************************************************************/
   AND_GATE #(.BubblesMask(2'b00))
      GATES_1 (.input1(s_logisimNet14),
               .input2(s_logisimNet23),
               .result(s_logisimNet15));

   OR_GATE_5_INPUTS #(.BubblesMask({1'b0, 4'h0}))
      GATES_2 (.input1(s_logisimNet6),
               .input2(s_logisimNet5),
               .input3(s_logisimNet2),
               .input4(s_logisimNet11),
               .input5(s_logisimNet18),
               .result(s_logisimNet17));

   Multiplexer_bus_2 #(.nrOfBits(32))
      PLEXERS_3 (.enable(1'b1),
                 .muxIn_0(s_logisimBus16[31:0]),
                 .muxIn_1(s_logisimBus12[31:0]),
                 .muxOut(s_logisimBus8[31:0]),
                 .sel(s_logisimNet6));

   Multiplexer_bus_2 #(.nrOfBits(32))
      PLEXERS_4 (.enable(1'b1),
                 .muxIn_0(s_logisimBus0[31:0]),
                 .muxIn_1(s_logisimBus8[31:0]),
                 .muxOut(s_logisimBus19[31:0]),
                 .sel(s_logisimNet17));

   Multiplexer_bus_2 #(.nrOfBits(32))
      PLEXERS_5 (.enable(1'b1),
                 .muxIn_0(s_logisimBus19[31:0]),
                 .muxIn_1(s_logisimBus20[31:0]),
                 .muxOut(s_logisimBus3[31:0]),
                 .sel(s_logisimNet21));

   Subtractor #(.extendedBits(33),
                .nrOfBits(32))
      ARITH_6 (.borrowIn(1'b0),
               .borrowOut(),
               .dataA(s_logisimBus9[31:0]),
               .dataB(s_logisimBus29[31:0]),
               .result(s_logisimBus4[31:0]));

   Comparator #(.nrOfBits(32),
                .twosComplement(1))
      ARITH_7 (.aEqualsB(s_logisimNet7),
               .aGreaterThanB(),
               .aLessThanB(),
               .dataA(s_logisimBus0[31:0]),
               .dataB(s_logisimBus10[31:0]));

   Comparator #(.nrOfBits(32),
                .twosComplement(1))
      ARITH_8 (.aEqualsB(s_logisimNet23),
               .aGreaterThanB(),
               .aLessThanB(),
               .dataA(s_logisimBus3[31:0]),
               .dataB(s_logisimBus10[31:0]));

   Comparator #(.nrOfBits(32),
                .twosComplement(1))
      ARITH_9 (.aEqualsB(),
               .aGreaterThanB(s_logisimNet21),
               .aLessThanB(),
               .dataA(s_logisimBus9[31:0]),
               .dataB(s_logisimBus1[31:0]));

   Shifter_32_bit #(.shifterMode(2))
      ARITH_10 (.dataA(s_logisimBus0[31:0]),
                .result(s_logisimBus13[31:0]),
                .shiftAmount(s_logisimBus22[4:0]));

   Shifter_32_bit #(.shifterMode(2))
      ARITH_11 (.dataA(s_logisimBus0[31:0]),
                .result(s_logisimBus12[31:0]),
                .shiftAmount(s_logisimBus30[4:0]));

   Shifter_32_bit #(.shifterMode(2))
      ARITH_12 (.dataA(s_logisimBus13[31:0]),
                .result(s_logisimBus16[31:0]),
                .shiftAmount(s_logisimBus31[4:0]));


endmodule
