/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
aluop
**
**
**
*****************************************************************************/
module
aluop(
Itype,
func,
op
);
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
Itype;
input
[5:0]
func;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
[3:0]
op;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
[3:0]
s_logisimBus0;
wire
[5:0]
s_logisimBus1;
wire
[3:0]
s_logisimBus10;
wire
[3:0]
s_logisimBus11;
wire
[3:0]
s_logisimBus12;
wire
[3:0]
s_logisimBus15;
wire
[3:0]
s_logisimBus17;
wire
[3:0]
s_logisimBus18;
wire
[3:0]
s_logisimBus19;
wire
[3:0]
s_logisimBus20;
wire
[3:0]
s_logisimBus21;
wire
[3:0]
s_logisimBus22;
wire
[3:0]
s_logisimBus23;
wire
[3:0]
s_logisimBus24;
wire
[3:0]
s_logisimBus25;
wire
[5:0]
s_logisimBus26;
wire
[5:0]
s_logisimBus27;
wire
[5:0]
s_logisimBus28;
wire
[5:0]
s_logisimBus29;
wire
[5:0]
s_logisimBus30;
wire
[5:0]
s_logisimBus31;
wire
[5:0]
s_logisimBus32;
wire
[5:0]
s_logisimBus33;
wire
[3:0]
s_logisimBus6;
wire
[3:0]
s_logisimBus8;
wire
[3:0]
s_logisimBus9;
wire
s_logisimNet13;
wire
s_logisimNet14;
wire
s_logisimNet16;
wire
s_logisimNet2;
wire
s_logisimNet3;
wire
s_logisimNet4;
wire
s_logisimNet5;
wire
s_logisimNet7;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
all
input
connections
are
defined
**
*******************************************************************************/
assign
s_logisimBus1[5:0]
=
func;
assign
s_logisimNet5
=
Itype;
/*******************************************************************************
**
Here
all
output
connections
are
defined
**
*******************************************************************************/
assign
op
=
s_logisimBus0[3:0];
/*******************************************************************************
**
Here
all
in-lined
components
are
defined
**
*******************************************************************************/
assign
s_logisimBus26[5:0]
=
{2'b10,
4'h2};
assign
s_logisimBus27[5:0]
=
{2'b10,
4'h4};
assign
s_logisimBus28[5:0]
=
{2'b10,
4'h5};
assign
s_logisimBus29[5:0]
=
{2'b10,
4'h6};
assign
s_logisimBus30[5:0]
=
{2'b00,
4'h4};
assign
s_logisimBus31[5:0]
=
{2'b00,
4'h6};
assign
s_logisimBus32[5:0]
=
{2'b00,
4'h7};
assign
s_logisimBus33[5:0]
=
{2'b10,
4'h0};
assign
s_logisimBus17[3:0]
=
4'h0;
assign
s_logisimBus18[3:0]
=
4'h1;
assign
s_logisimBus19[3:0]
=
4'h4;
assign
s_logisimBus20[3:0]
=
4'h5;
assign
s_logisimBus21[3:0]
=
4'h6;
assign
s_logisimBus22[3:0]
=
4'h9;
assign
s_logisimBus23[3:0]
=
4'hA;
assign
s_logisimBus24[3:0]
=
4'hB;
assign
s_logisimBus25[3:0]
=
4'hC;
/*******************************************************************************
**
Here
all
normal
components
are
defined
**
*******************************************************************************/
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_1
(.enable(1'b1),
.muxIn_0(s_logisimBus17[3:0]),
.muxIn_1(s_logisimBus18[3:0]),
.muxOut(s_logisimBus12[3:0]),
.sel(s_logisimNet13));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_2
(.enable(1'b1),
.muxIn_0(s_logisimBus12[3:0]),
.muxIn_1(s_logisimBus19[3:0]),
.muxOut(s_logisimBus8[3:0]),
.sel(s_logisimNet3));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_3
(.enable(1'b1),
.muxIn_0(s_logisimBus8[3:0]),
.muxIn_1(s_logisimBus20[3:0]),
.muxOut(s_logisimBus9[3:0]),
.sel(s_logisimNet7));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_4
(.enable(1'b1),
.muxIn_0(s_logisimBus9[3:0]),
.muxIn_1(s_logisimBus21[3:0]),
.muxOut(s_logisimBus10[3:0]),
.sel(s_logisimNet2));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_5
(.enable(1'b1),
.muxIn_0(s_logisimBus10[3:0]),
.muxIn_1(s_logisimBus22[3:0]),
.muxOut(s_logisimBus11[3:0]),
.sel(s_logisimNet16));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_6
(.enable(1'b1),
.muxIn_0(s_logisimBus11[3:0]),
.muxIn_1(s_logisimBus23[3:0]),
.muxOut(s_logisimBus15[3:0]),
.sel(s_logisimNet4));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_7
(.enable(1'b1),
.muxIn_0(s_logisimBus15[3:0]),
.muxIn_1(s_logisimBus24[3:0]),
.muxOut(s_logisimBus6[3:0]),
.sel(s_logisimNet14));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_8
(.enable(1'b1),
.muxIn_0(s_logisimBus6[3:0]),
.muxIn_1(s_logisimBus25[3:0]),
.muxOut(s_logisimBus0[3:0]),
.sel(s_logisimNet5));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_9
(.aEqualsB(s_logisimNet13),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus26[5:0]),
.dataB(s_logisimBus1[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_10
(.aEqualsB(s_logisimNet3),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus27[5:0]),
.dataB(s_logisimBus1[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_11
(.aEqualsB(s_logisimNet7),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus28[5:0]),
.dataB(s_logisimBus1[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_12
(.aEqualsB(s_logisimNet2),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus29[5:0]),
.dataB(s_logisimBus1[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_13
(.aEqualsB(s_logisimNet16),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus30[5:0]),
.dataB(s_logisimBus1[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_14
(.aEqualsB(s_logisimNet4),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus31[5:0]),
.dataB(s_logisimBus1[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_15
(.aEqualsB(s_logisimNet14),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus32[5:0]),
.dataB(s_logisimBus1[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_16
(.aEqualsB(),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus33[5:0]),
.dataB(s_logisimBus1[5:0]));
endmodule