/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
BitSelector
**
**
**
*****************************************************************************/
module
BitSelector(
dataIn,
dataOut,
sel
);
/*******************************************************************************
**
Here
all
module
parameters
are
defined
with
a
dummy
value
**
*******************************************************************************/
parameter
nrOfExtendedBits
=
1;
parameter
nrOfInputBits
=
1;
parameter
nrOfselBits
=
1;
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
[nrOfInputBits-1:0]
dataIn;
input
[nrOfselBits-1:0]
sel;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
dataOut;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
[nrOfExtendedBits-1:0]
s_extendedVector;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
assign
s_extendedVector[nrOfExtendedBits-1:nrOfInputBits]
=
0;
assign
s_extendedVector[nrOfInputBits-1:0]
=
dataIn;
assign
dataOut
=
s_extendedVector[sel];
endmodule