/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
find_msb
**
**
**
*****************************************************************************/
module
find_msb(
input1,
result_msb
);
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
[63:0]
input1;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
[7:0]
result_msb;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
[5:0]
s_logisimBus1;
wire
[5:0]
s_logisimBus100;
wire
[5:0]
s_logisimBus101;
wire
[5:0]
s_logisimBus102;
wire
[5:0]
s_logisimBus103;
wire
[5:0]
s_logisimBus104;
wire
[5:0]
s_logisimBus106;
wire
[5:0]
s_logisimBus108;
wire
[5:0]
s_logisimBus109;
wire
[5:0]
s_logisimBus11;
wire
[5:0]
s_logisimBus110;
wire
[5:0]
s_logisimBus111;
wire
[5:0]
s_logisimBus112;
wire
[5:0]
s_logisimBus113;
wire
[5:0]
s_logisimBus114;
wire
[5:0]
s_logisimBus115;
wire
[5:0]
s_logisimBus116;
wire
[5:0]
s_logisimBus118;
wire
[5:0]
s_logisimBus119;
wire
[5:0]
s_logisimBus12;
wire
[5:0]
s_logisimBus120;
wire
[5:0]
s_logisimBus121;
wire
[5:0]
s_logisimBus122;
wire
[5:0]
s_logisimBus123;
wire
[5:0]
s_logisimBus128;
wire
[5:0]
s_logisimBus13;
wire
[5:0]
s_logisimBus130;
wire
[5:0]
s_logisimBus131;
wire
[5:0]
s_logisimBus133;
wire
[5:0]
s_logisimBus134;
wire
[5:0]
s_logisimBus135;
wire
[5:0]
s_logisimBus137;
wire
[5:0]
s_logisimBus138;
wire
[5:0]
s_logisimBus139;
wire
[5:0]
s_logisimBus140;
wire
[5:0]
s_logisimBus142;
wire
[5:0]
s_logisimBus143;
wire
[5:0]
s_logisimBus144;
wire
[5:0]
s_logisimBus145;
wire
[5:0]
s_logisimBus146;
wire
[5:0]
s_logisimBus147;
wire
[5:0]
s_logisimBus148;
wire
[5:0]
s_logisimBus150;
wire
[5:0]
s_logisimBus151;
wire
[5:0]
s_logisimBus152;
wire
[5:0]
s_logisimBus153;
wire
[5:0]
s_logisimBus155;
wire
[5:0]
s_logisimBus156;
wire
[5:0]
s_logisimBus158;
wire
[5:0]
s_logisimBus159;
wire
[5:0]
s_logisimBus16;
wire
[5:0]
s_logisimBus160;
wire
[5:0]
s_logisimBus161;
wire
[5:0]
s_logisimBus163;
wire
[5:0]
s_logisimBus164;
wire
[5:0]
s_logisimBus166;
wire
[5:0]
s_logisimBus168;
wire
[5:0]
s_logisimBus17;
wire
[5:0]
s_logisimBus170;
wire
[5:0]
s_logisimBus171;
wire
[5:0]
s_logisimBus172;
wire
[5:0]
s_logisimBus173;
wire
[5:0]
s_logisimBus175;
wire
[5:0]
s_logisimBus177;
wire
[5:0]
s_logisimBus178;
wire
[5:0]
s_logisimBus18;
wire
[5:0]
s_logisimBus181;
wire
[5:0]
s_logisimBus182;
wire
[5:0]
s_logisimBus183;
wire
[5:0]
s_logisimBus184;
wire
[5:0]
s_logisimBus185;
wire
[63:0]
s_logisimBus187;
wire
[5:0]
s_logisimBus188;
wire
[5:0]
s_logisimBus189;
wire
[5:0]
s_logisimBus19;
wire
[5:0]
s_logisimBus190;
wire
[5:0]
s_logisimBus191;
wire
[5:0]
s_logisimBus192;
wire
[5:0]
s_logisimBus193;
wire
[5:0]
s_logisimBus194;
wire
[5:0]
s_logisimBus195;
wire
[5:0]
s_logisimBus2;
wire
[5:0]
s_logisimBus20;
wire
[5:0]
s_logisimBus21;
wire
[5:0]
s_logisimBus22;
wire
[5:0]
s_logisimBus23;
wire
[5:0]
s_logisimBus24;
wire
[5:0]
s_logisimBus25;
wire
[5:0]
s_logisimBus26;
wire
[5:0]
s_logisimBus27;
wire
[5:0]
s_logisimBus28;
wire
[5:0]
s_logisimBus29;
wire
[5:0]
s_logisimBus3;
wire
[5:0]
s_logisimBus34;
wire
[5:0]
s_logisimBus35;
wire
[5:0]
s_logisimBus36;
wire
[5:0]
s_logisimBus39;
wire
[5:0]
s_logisimBus4;
wire
[5:0]
s_logisimBus40;
wire
[5:0]
s_logisimBus41;
wire
[5:0]
s_logisimBus42;
wire
[5:0]
s_logisimBus43;
wire
[5:0]
s_logisimBus45;
wire
[5:0]
s_logisimBus46;
wire
[5:0]
s_logisimBus47;
wire
[5:0]
s_logisimBus48;
wire
[5:0]
s_logisimBus49;
wire
[5:0]
s_logisimBus50;
wire
[5:0]
s_logisimBus51;
wire
[5:0]
s_logisimBus52;
wire
[5:0]
s_logisimBus53;
wire
[5:0]
s_logisimBus55;
wire
[5:0]
s_logisimBus57;
wire
[5:0]
s_logisimBus58;
wire
[5:0]
s_logisimBus6;
wire
[5:0]
s_logisimBus60;
wire
[5:0]
s_logisimBus62;
wire
[5:0]
s_logisimBus64;
wire
[5:0]
s_logisimBus65;
wire
[5:0]
s_logisimBus67;
wire
[5:0]
s_logisimBus68;
wire
[5:0]
s_logisimBus69;
wire
[5:0]
s_logisimBus7;
wire
[5:0]
s_logisimBus70;
wire
[7:0]
s_logisimBus72;
wire
[5:0]
s_logisimBus73;
wire
[5:0]
s_logisimBus74;
wire
[5:0]
s_logisimBus75;
wire
[7:0]
s_logisimBus76;
wire
[5:0]
s_logisimBus77;
wire
[5:0]
s_logisimBus78;
wire
[5:0]
s_logisimBus79;
wire
[7:0]
s_logisimBus8;
wire
[5:0]
s_logisimBus82;
wire
[5:0]
s_logisimBus84;
wire
[5:0]
s_logisimBus86;
wire
[5:0]
s_logisimBus87;
wire
[5:0]
s_logisimBus88;
wire
[5:0]
s_logisimBus9;
wire
[5:0]
s_logisimBus90;
wire
[5:0]
s_logisimBus91;
wire
[5:0]
s_logisimBus92;
wire
[5:0]
s_logisimBus93;
wire
[5:0]
s_logisimBus94;
wire
[5:0]
s_logisimBus95;
wire
[5:0]
s_logisimBus97;
wire
s_logisimNet0;
wire
s_logisimNet10;
wire
s_logisimNet105;
wire
s_logisimNet107;
wire
s_logisimNet117;
wire
s_logisimNet124;
wire
s_logisimNet125;
wire
s_logisimNet126;
wire
s_logisimNet127;
wire
s_logisimNet129;
wire
s_logisimNet132;
wire
s_logisimNet136;
wire
s_logisimNet14;
wire
s_logisimNet141;
wire
s_logisimNet149;
wire
s_logisimNet15;
wire
s_logisimNet154;
wire
s_logisimNet157;
wire
s_logisimNet162;
wire
s_logisimNet165;
wire
s_logisimNet167;
wire
s_logisimNet169;
wire
s_logisimNet174;
wire
s_logisimNet176;
wire
s_logisimNet179;
wire
s_logisimNet180;
wire
s_logisimNet186;
wire
s_logisimNet30;
wire
s_logisimNet31;
wire
s_logisimNet32;
wire
s_logisimNet33;
wire
s_logisimNet37;
wire
s_logisimNet38;
wire
s_logisimNet44;
wire
s_logisimNet5;
wire
s_logisimNet56;
wire
s_logisimNet59;
wire
s_logisimNet61;
wire
s_logisimNet63;
wire
s_logisimNet71;
wire
s_logisimNet80;
wire
s_logisimNet81;
wire
s_logisimNet83;
wire
s_logisimNet85;
wire
s_logisimNet89;
wire
s_logisimNet96;
wire
s_logisimNet98;
wire
s_logisimNet99;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
all
input
connections
are
defined
**
*******************************************************************************/
assign
s_logisimBus187[63:0]
=
input1;
/*******************************************************************************
**
Here
all
output
connections
are
defined
**
*******************************************************************************/
assign
result_msb
=
s_logisimBus8[7:0];
/*******************************************************************************
**
Here
all
in-lined
components
are
defined
**
*******************************************************************************/
assign
s_logisimBus158[5:0]
=
{2'b10,
4'h6};
assign
s_logisimBus182[5:0]
=
{2'b00,
4'h8};
assign
s_logisimBus121[5:0]
=
{2'b10,
4'h5};
assign
s_logisimBus148[5:0]
=
{2'b00,
4'h9};
assign
s_logisimBus78[5:0]
=
{2'b10,
4'h4};
assign
s_logisimBus102[5:0]
=
{2'b00,
4'hA};
assign
s_logisimBus24[5:0]
=
{2'b10,
4'h3};
assign
s_logisimBus52[5:0]
=
{2'b00,
4'hB};
assign
s_logisimBus168[5:0]
=
{2'b10,
4'h2};
assign
s_logisimBus193[5:0]
=
{2'b00,
4'hC};
assign
s_logisimBus118[5:0]
=
{2'b10,
4'h1};
assign
s_logisimBus146[5:0]
=
{2'b00,
4'hD};
assign
s_logisimBus116[5:0]
=
{2'b10,
4'h0};
assign
s_logisimBus142[5:0]
=
{2'b00,
4'hE};
assign
s_logisimBus93[5:0]
=
{2'b11,
4'hE};
assign
s_logisimBus139[5:0]
=
{2'b10,
4'hE};
assign
s_logisimBus164[5:0]
=
{2'b00,
4'h0};
assign
s_logisimBus143[5:0]
=
{2'b01,
4'hF};
assign
s_logisimBus166[5:0]
=
{2'b00,
4'hF};
assign
s_logisimBus23[5:0]
=
{2'b01,
4'hE};
assign
s_logisimBus48[5:0]
=
{2'b01,
4'h0};
assign
s_logisimBus94[5:0]
=
{2'b01,
4'hD};
assign
s_logisimBus115[5:0]
=
{2'b01,
4'h1};
assign
s_logisimBus50[5:0]
=
{2'b01,
4'hC};
assign
s_logisimBus73[5:0]
=
{2'b01,
4'h2};
assign
s_logisimBus175[5:0]
=
{2'b01,
4'hB};
assign
s_logisimBus3[5:0]
=
{2'b01,
4'h3};
assign
s_logisimBus4[5:0]
=
{2'b01,
4'hA};
assign
s_logisimBus34[5:0]
=
{2'b01,
4'h4};
assign
s_logisimBus150[5:0]
=
{2'b01,
4'h9};
assign
s_logisimBus171[5:0]
=
{2'b01,
4'h5};
assign
s_logisimBus151[5:0]
=
{2'b01,
4'h8};
assign
s_logisimBus172[5:0]
=
{2'b01,
4'h6};
assign
s_logisimBus152[5:0]
=
{2'b01,
4'h7};
assign
s_logisimBus173[5:0]
=
{2'b01,
4'h7};
assign
s_logisimBus29[5:0]
=
{2'b01,
4'h6};
assign
s_logisimBus57[5:0]
=
{2'b01,
4'h8};
assign
s_logisimBus20[5:0]
=
{2'b10,
4'hD};
assign
s_logisimBus45[5:0]
=
{2'b00,
4'h1};
assign
s_logisimBus170[5:0]
=
{2'b01,
4'h5};
assign
s_logisimBus2[5:0]
=
{2'b01,
4'h9};
assign
s_logisimBus1[5:0]
=
{2'b01,
4'h4};
assign
s_logisimBus26[5:0]
=
{2'b01,
4'hA};
assign
s_logisimBus27[5:0]
=
{2'b01,
4'h3};
assign
s_logisimBus55[5:0]
=
{2'b01,
4'hB};
assign
s_logisimBus130[5:0]
=
{2'b01,
4'h2};
assign
s_logisimBus155[5:0]
=
{2'b01,
4'hC};
assign
s_logisimBus40[5:0]
=
{2'b01,
4'h1};
assign
s_logisimBus64[5:0]
=
{2'b01,
4'hD};
assign
s_logisimBus60[5:0]
=
{2'b01,
4'h0};
assign
s_logisimBus84[5:0]
=
{2'b01,
4'hE};
assign
s_logisimBus13[5:0]
=
{2'b00,
4'hF};
assign
s_logisimBus39[5:0]
=
{2'b01,
4'hF};
assign
s_logisimBus101[5:0]
=
{2'b00,
4'hE};
assign
s_logisimBus122[5:0]
=
{2'b10,
4'h0};
assign
s_logisimBus161[5:0]
=
{2'b10,
4'hC};
assign
s_logisimBus185[5:0]
=
{2'b00,
4'h2};
assign
s_logisimBus153[5:0]
=
{2'b00,
4'hD};
assign
s_logisimBus178[5:0]
=
{2'b10,
4'h1};
assign
s_logisimBus7[5:0]
=
{2'b00,
4'hC};
assign
s_logisimBus35[5:0]
=
{2'b10,
4'h2};
assign
s_logisimBus36[5:0]
=
{2'b00,
4'hB};
assign
s_logisimBus58[5:0]
=
{2'b10,
4'h3};
assign
s_logisimBus47[5:0]
=
{2'b00,
4'hA};
assign
s_logisimBus22[5:0]
=
{2'b10,
4'h4};
assign
s_logisimBus140[5:0]
=
{2'b00,
4'h9};
assign
s_logisimBus113[5:0]
=
{2'b10,
4'h5};
assign
s_logisimBus184[5:0]
=
{2'b00,
4'h8};
assign
s_logisimBus160[5:0]
=
{2'b10,
4'h6};
assign
s_logisimBus21[5:0]
=
{2'b00,
4'h7};
assign
s_logisimBus92[5:0]
=
{2'b10,
4'h7};
assign
s_logisimBus137[5:0]
=
{2'b00,
4'h6};
assign
s_logisimBus111[5:0]
=
{2'b10,
4'h8};
assign
s_logisimBus90[5:0]
=
{2'b00,
4'h5};
assign
s_logisimBus65[5:0]
=
{2'b10,
4'h9};
assign
s_logisimBus112[5:0]
=
{2'b10,
4'hB};
assign
s_logisimBus138[5:0]
=
{2'b00,
4'h3};
assign
s_logisimBus68[5:0]
=
{2'b00,
4'h4};
assign
s_logisimBus134[5:0]
=
{2'b10,
4'hA};
assign
s_logisimBus17[5:0]
=
{2'b00,
4'h3};
assign
s_logisimBus86[5:0]
=
{2'b10,
4'hB};
assign
s_logisimBus42[5:0]
=
{2'b00,
4'h2};
assign
s_logisimBus19[5:0]
=
{2'b10,
4'hC};
assign
s_logisimBus147[5:0]
=
{2'b00,
4'h1};
assign
s_logisimBus120[5:0]
=
{2'b10,
4'hD};
assign
s_logisimBus123[5:0]
=
{2'b00,
4'h0};
assign
s_logisimBus194[5:0]
=
{2'b10,
4'hE};
assign
s_logisimBus72[7:6]
=
2'b00;
assign
s_logisimBus76[7:0]
=
8'hFF;
assign
s_logisimBus145[5:0]
=
{2'b10,
4'hF};
assign
s_logisimBus67[5:0]
=
{2'b10,
4'hA};
assign
s_logisimBus91[5:0]
=
{2'b00,
4'h4};
assign
s_logisimBus135[5:0]
=
{2'b10,
4'h9};
assign
s_logisimBus159[5:0]
=
{2'b00,
4'h5};
assign
s_logisimBus87[5:0]
=
{2'b10,
4'h8};
assign
s_logisimBus108[5:0]
=
{2'b00,
4'h6};
assign
s_logisimBus18[5:0]
=
{2'b10,
4'h7};
assign
s_logisimBus41[5:0]
=
{2'b00,
4'h7};
/*******************************************************************************
**
Here
all
normal
components
are
defined
**
*******************************************************************************/
BitSelector
#(.nrOfExtendedBits(65),
.nrOfInputBits(64),
.nrOfselBits(6))
PLEXERS_1
(.dataIn(s_logisimBus187[63:0]),
.dataOut(s_logisimNet83),
.sel(s_logisimBus182[5:0]));
Multiplexer_bus_2
#(.nrOfBits(6))
PLEXERS_2
(.enable(1'b1),
.muxIn_0(s_logisimBus195[5:0]),
.muxIn_1(s_logisimBus158[5:0]),
.muxOut(s_logisimBus131[5:0]),
.sel(s_logisimNet83));
BitSelector
#(.nrOfExtendedBits(65),
.nrOfInputBits(64),
.nrOfselBits(6))
PLEXERS_3
(.dataIn(s_logisimBus187[63:0]),
.dataOut(s_logisimNet33),
.sel(s_logisimBus148[5:0]));
Multiplexer_bus_2
#(.nrOfBits(6))
PLEXERS_4
(.enable(1'b1),
.muxIn_0(s_logisimBus131[5:0]),
.muxIn_1(s_logisimBus121[5:0]),
.muxOut(s_logisimBus88[5:0]),
.sel(s_logisimNet33));
BitSelector
#(.nrOfExtendedBits(65),
.nrOfInputBits(64),
.nrOfselBits(6))
PLEXERS_5
(.dataIn(s_logisimBus187[63:0]),
.dataOut(s_logisimNet174),
.sel(s_logisimBus102[5:0]));
Multiplexer_bus_2
#(.nrOfBits(6))
PLEXERS_6
(.enable(1'b1),
.muxIn_0(s_logisimBus88[5:0]),
.muxIn_1(s_logisimBus78[5:0]),
.muxOut(s_logisimBus43[5:0]),
.sel(s_logisimNet174));
BitSelector
#(.nrOfExtendedBits(65),
.nrOfInputBits(64),
.nrOfselBits(6))
PLEXERS_7
(.dataIn(s_logisimBus187[63:0]),
.dataOut(s_logisimNet126),
.sel(s_logisimBus52[5:0]));
Multiplexer_bus_2
#(.nrOfBits(6))
PLEXERS_8
(.enable(1'b1),
.muxIn_0(s_logisimBus43[5:0]),
.muxIn_1(s_logisimBus24[5:0]),
.muxOut(s_logisimBus183[5:0]),
.sel(s_logisimNet126));
BitSelector
#(.nrOfExtendedBits(65),
.nrOfInputBits(64),
.nrOfselBits(6))
PLEXERS_9
(.dataIn(s_logisimBus187[63:0]),
.dataOut(s_logisimNet80),
.sel(s_logisimBus193[5:0]));
Multiplexer_bus_2
#(.nrOfBits(6))
PLEXERS_10
(.enable(1'b1),
.muxIn_0(s_logisimBus183[5:0]),
.muxIn_1(s_logisimBus168[5:0]),
.muxOut(s_logisimBus133[5:0]),
.sel(s_logisimNet80));
BitSelector
#(.nrOfExtendedBits(65),
.nrOfInputBits(64),
.nrOfselBits(6))
PLEXERS_11
(.dataIn(s_logisimBus187[63:0]),
.dataOut(s_logisimNet30),
.sel(s_logisimBus146[5:0]));
Multiplexer_bus_2
#(.nrOfBits(6))
PLEXERS_12
(.enable(1'b1),
.muxIn_0(s_logisimBus133[5:0]),
.muxIn_1(s_logisimBus118[5:0]),
.muxOut(s_logisimBus62[5:0]),
.sel(s_logisimNet30));
BitSelector
#(.nrOfExtendedBits(65),
.nrOfInputBits(64),
.nrOfselBits(6))
PLEXERS_13
(.dataIn(s_logisimBus187[63:0]),
.dataOut(s_logisimNet31),
.sel(s_logisimBus142[5:0]));
Multiplexer_bus_2
#(.nrOfBits(6))
PLEXERS_14
(.enable(1'b1),
.muxIn_0(s_logisimBus62[5:0]),
.muxIn_1(s_logisimBus116[5:0]),
.muxOut(s_logisimBus25[5:0]),
.sel(s_logisimNet31));
BitSelector
#(.nrOfExtendedBits(65),
.nrOfInputBits(64),
.nrOfselBits(6))
PLEXERS_15
(.dataIn(s_logisimBus187[63:0]),
.dataOut(s_logisimNet56),
.sel(s_logisimBus166[5:0]));
Multiplexer_bus_2
#(.nrOfBits(6))
PLEXERS_16
(.enable(1'b1),
.muxIn_0(s_logisimBus25[5:0]),
.muxIn_1(s_logisimBus143[5:0]),
.muxOut(s_logisimBus181[5:0]),
.sel(s_logisimNet56));
BitSelector
#(.nrOfExtendedBits(65),
.nrOfInputBits(64),
.nrOfselBits(6))
PLEXERS_17
(.dataIn(s_logisimBus187[63:0]),
.dataOut(s_logisimNet125),
.sel(s_logisimBus48[5:0]));
Multiplexer_bus_2
#(.nrOfBits(6))
PLEXERS_18
(.enable(1'b1),
.muxIn_0(s_logisimBus181[5:0]),
.muxIn_1(s_logisimBus23[5:0]),
.muxOut(s_logisimBus69[5:0]),
.sel(s_logisimNet125));
BitSelector
#(.nrOfExtendedBits(65),
.nrOfInputBits(64),
.nrOfselBits(6))
PLEXERS_19
(.dataIn(s_logisimBus187[63:0]),
.dataOut(s_logisimNet0),
.sel(s_logisimBus115[5:0]));
BitSelector
#(.nrOfExtendedBits(65),
.nrOfInputBits(64),
.nrOfselBits(6))
PLEXERS_20
(.dataIn(s_logisimBus187[63:0]),
.dataOut(s_logisimNet63),
.sel(s_logisimBus164[5:0]));
Multiplexer_bus_2
#(.nrOfBits(6))
PLEXERS_21
(.enable(1'b1),
.muxIn_0(s_logisimBus69[5:0]),
.muxIn_1(s_logisimBus94[5:0]),
.muxOut(s_logisimBus70[5:0]),
.sel(s_logisimNet0));
BitSelector
#(.nrOfExtendedBits(65),
.nrOfInputBits(64),
.nrOfselBits(6))
PLEXERS_22
(.dataIn(s_logisimBus187[63:0]),
.dataOut(s_logisimNet169),
.sel(s_logisimBus73[5:0]));
Multiplexer_bus_2
#(.nrOfBits(6))
PLEXERS_23
(.enable(1'b1),
.muxIn_0(s_logisimBus70[5:0]),
.muxIn_1(s_logisimBus50[5:0]),
.muxOut(s_logisimBus6[5:0]),
.sel(s_logisimNet169));
Multiplexer_bus_2
#(.nrOfBits(6))
PLEXERS_24
(.enable(1'b1),
.muxIn_0(s_logisimBus93[5:0]),
.muxIn_1(s_logisimBus139[5:0]),
.muxOut(s_logisimBus192[5:0]),
.sel(s_logisimNet63));
BitSelector
#(.nrOfExtendedBits(65),
.nrOfInputBits(64),
.nrOfselBits(6))
PLEXERS_25
(.dataIn(s_logisimBus187[63:0]),
.dataOut(s_logisimNet124),
.sel(s_logisimBus3[5:0]));
Multiplexer_bus_2
#(.nrOfBits(6))
PLEXERS_26
(.enable(1'b1),
.muxIn_0(s_logisimBus6[5:0]),
.muxIn_1(s_logisimBus175[5:0]),
.muxOut(s_logisimBus79[5:0]),
.sel(s_logisimNet124));
BitSelector
#(.nrOfExtendedBits(65),
.nrOfInputBits(64),
.nrOfselBits(6))
PLEXERS_27
(.dataIn(s_logisimBus187[63:0]),
.dataOut(s_logisimNet149),
.sel(s_logisimBus34[5:0]));
Multiplexer_bus_2
#(.nrOfBits(6))
PLEXERS_28
(.enable(1'b1),
.muxIn_0(s_logisimBus79[5:0]),
.muxIn_1(s_logisimBus4[5:0]),
.muxOut(s_logisimBus177[5:0]),
.sel(s_logisimNet149));
BitSelector
#(.nrOfExtendedBits(65),
.nrOfInputBits(64),
.nrOfselBits(6))
PLEXERS_29
(.dataIn(s_logisimBus187[63:0]),
.dataOut(s_logisimNet99),
.sel(s_logisimBus171[5:0]));
Multiplexer_bus_2
#(.nrOfBits(6))
PLEXERS_30
(.enable(1'b1),
.muxIn_0(s_logisimBus177[5:0]),
.muxIn_1(s_logisimBus150[5:0]),
.muxOut(s_logisimBus109[5:0]),
.sel(s_logisimNet99));
BitSelector
#(.nrOfExtendedBits(65),
.nrOfInputBits(64),
.nrOfselBits(6))
PLEXERS_31
(.dataIn(s_logisimBus187[63:0]),
.dataOut(s_logisimNet96),
.sel(s_logisimBus172[5:0]));
Multiplexer_bus_2
#(.nrOfBits(6))
PLEXERS_32
(.enable(1'b1),
.muxIn_0(s_logisimBus109[5:0]),
.muxIn_1(s_logisimBus151[5:0]),
.muxOut(s_logisimBus110[5:0]),
.sel(s_logisimNet96));
BitSelector
#(.nrOfExtendedBits(65),
.nrOfInputBits(64),
.nrOfselBits(6))
PLEXERS_33
(.dataIn(s_logisimBus187[63:0]),
.dataOut(s_logisimNet98),
.sel(s_logisimBus173[5:0]));
Multiplexer_bus_2
#(.nrOfBits(6))
PLEXERS_34
(.enable(1'b1),
.muxIn_0(s_logisimBus110[5:0]),
.muxIn_1(s_logisimBus152[5:0]),
.muxOut(s_logisimBus9[5:0]),
.sel(s_logisimNet98));
BitSelector
#(.nrOfExtendedBits(65),
.nrOfInputBits(64),
.nrOfselBits(6))
PLEXERS_35
(.dataIn(s_logisimBus187[63:0]),
.dataOut(s_logisimNet167),
.sel(s_logisimBus57[5:0]));
Multiplexer_bus_2
#(.nrOfBits(6))
PLEXERS_36
(.enable(1'b1),
.muxIn_0(s_logisimBus9[5:0]),
.muxIn_1(s_logisimBus29[5:0]),
.muxOut(s_logisimBus12[5:0]),
.sel(s_logisimNet167));
BitSelector
#(.nrOfExtendedBits(65),
.nrOfInputBits(64),
.nrOfselBits(6))
PLEXERS_37
(.dataIn(s_logisimBus187[63:0]),
.dataOut(s_logisimNet117),
.sel(s_logisimBus2[5:0]));
Multiplexer_bus_2
#(.nrOfBits(6))
PLEXERS_38
(.enable(1'b1),
.muxIn_0(s_logisimBus12[5:0]),
.muxIn_1(s_logisimBus170[5:0]),
.muxOut(s_logisimBus82[5:0]),
.sel(s_logisimNet117));
BitSelector
#(.nrOfExtendedBits(65),
.nrOfInputBits(64),
.nrOfselBits(6))
PLEXERS_39
(.dataIn(s_logisimBus187[63:0]),
.dataOut(s_logisimNet141),
.sel(s_logisimBus26[5:0]));
Multiplexer_bus_2
#(.nrOfBits(6))
PLEXERS_40
(.enable(1'b1),
.muxIn_0(s_logisimBus82[5:0]),
.muxIn_1(s_logisimBus1[5:0]),
.muxOut(s_logisimBus104[5:0]),
.sel(s_logisimNet141));
BitSelector
#(.nrOfExtendedBits(65),
.nrOfInputBits(64),
.nrOfselBits(6))
PLEXERS_41
(.dataIn(s_logisimBus187[63:0]),
.dataOut(s_logisimNet129),
.sel(s_logisimBus45[5:0]));
BitSelector
#(.nrOfExtendedBits(65),
.nrOfInputBits(64),
.nrOfselBits(6))
PLEXERS_42
(.dataIn(s_logisimBus187[63:0]),
.dataOut(s_logisimNet165),
.sel(s_logisimBus55[5:0]));
Multiplexer_bus_2
#(.nrOfBits(6))
PLEXERS_43
(.enable(1'b1),
.muxIn_0(s_logisimBus104[5:0]),
.muxIn_1(s_logisimBus27[5:0]),
.muxOut(s_logisimBus74[5:0]),
.sel(s_logisimNet165));
Multiplexer_bus_2
#(.nrOfBits(6))
PLEXERS_44
(.enable(1'b1),
.muxIn_0(s_logisimBus192[5:0]),
.muxIn_1(s_logisimBus20[5:0]),
.muxOut(s_logisimBus191[5:0]),
.sel(s_logisimNet129));
BitSelector
#(.nrOfExtendedBits(65),
.nrOfInputBits(64),
.nrOfselBits(6))
PLEXERS_45
(.dataIn(s_logisimBus187[63:0]),
.dataOut(s_logisimNet71),
.sel(s_logisimBus155[5:0]));
Multiplexer_bus_2
#(.nrOfBits(6))
PLEXERS_46
(.enable(1'b1),
.muxIn_0(s_logisimBus74[5:0]),
.muxIn_1(s_logisimBus130[5:0]),
.muxOut(s_logisimBus163[5:0]),
.sel(s_logisimNet71));
BitSelector
#(.nrOfExtendedBits(65),
.nrOfInputBits(64),
.nrOfselBits(6))
PLEXERS_47
(.dataIn(s_logisimBus187[63:0]),
.dataOut(s_logisimNet162),
.sel(s_logisimBus64[5:0]));
Multiplexer_bus_2
#(.nrOfBits(6))
PLEXERS_48
(.enable(1'b1),
.muxIn_0(s_logisimBus163[5:0]),
.muxIn_1(s_logisimBus40[5:0]),
.muxOut(s_logisimBus128[5:0]),
.sel(s_logisimNet162));
BitSelector
#(.nrOfExtendedBits(65),
.nrOfInputBits(64),
.nrOfselBits(6))
PLEXERS_49
(.dataIn(s_logisimBus187[63:0]),
.dataOut(s_logisimNet186),
.sel(s_logisimBus84[5:0]));
Multiplexer_bus_2
#(.nrOfBits(6))
PLEXERS_50
(.enable(1'b1),
.muxIn_0(s_logisimBus128[5:0]),
.muxIn_1(s_logisimBus60[5:0]),
.muxOut(s_logisimBus28[5:0]),
.sel(s_logisimNet186));
BitSelector
#(.nrOfExtendedBits(65),
.nrOfInputBits(64),
.nrOfselBits(6))
PLEXERS_51
(.dataIn(s_logisimBus187[63:0]),
.dataOut(s_logisimNet136),
.sel(s_logisimBus39[5:0]));
Multiplexer_bus_2
#(.nrOfBits(6))
PLEXERS_52
(.enable(1'b1),
.muxIn_0(s_logisimBus28[5:0]),
.muxIn_1(s_logisimBus13[5:0]),
.muxOut(s_logisimBus46[5:0]),
.sel(s_logisimNet136));
BitSelector
#(.nrOfExtendedBits(65),
.nrOfInputBits(64),
.nrOfselBits(6))
PLEXERS_53
(.dataIn(s_logisimBus187[63:0]),
.dataOut(s_logisimNet44),
.sel(s_logisimBus122[5:0]));
Multiplexer_bus_2
#(.nrOfBits(6))
PLEXERS_54
(.enable(1'b1),
.muxIn_0(s_logisimBus46[5:0]),
.muxIn_1(s_logisimBus101[5:0]),
.muxOut(s_logisimBus190[5:0]),
.sel(s_logisimNet44));
BitSelector
#(.nrOfExtendedBits(65),
.nrOfInputBits(64),
.nrOfselBits(6))
PLEXERS_55
(.dataIn(s_logisimBus187[63:0]),
.dataOut(s_logisimNet89),
.sel(s_logisimBus178[5:0]));
Multiplexer_bus_2
#(.nrOfBits(6))
PLEXERS_56
(.enable(1'b1),
.muxIn_0(s_logisimBus190[5:0]),
.muxIn_1(s_logisimBus153[5:0]),
.muxOut(s_logisimBus49[5:0]),
.sel(s_logisimNet89));
BitSelector
#(.nrOfExtendedBits(65),
.nrOfInputBits(64),
.nrOfselBits(6))
PLEXERS_57
(.dataIn(s_logisimBus187[63:0]),
.dataOut(s_logisimNet132),
.sel(s_logisimBus35[5:0]));
Multiplexer_bus_2
#(.nrOfBits(6))
PLEXERS_58
(.enable(1'b1),
.muxIn_0(s_logisimBus49[5:0]),
.muxIn_1(s_logisimBus7[5:0]),
.muxOut(s_logisimBus106[5:0]),
.sel(s_logisimNet132));
BitSelector
#(.nrOfExtendedBits(65),
.nrOfInputBits(64),
.nrOfselBits(6))
PLEXERS_59
(.dataIn(s_logisimBus187[63:0]),
.dataOut(s_logisimNet85),
.sel(s_logisimBus185[5:0]));
BitSelector
#(.nrOfExtendedBits(65),
.nrOfInputBits(64),
.nrOfselBits(6))
PLEXERS_60
(.dataIn(s_logisimBus187[63:0]),
.dataOut(s_logisimNet157),
.sel(s_logisimBus58[5:0]));
Multiplexer_bus_2
#(.nrOfBits(6))
PLEXERS_61
(.enable(1'b1),
.muxIn_0(s_logisimBus106[5:0]),
.muxIn_1(s_logisimBus36[5:0]),
.muxOut(s_logisimBus188[5:0]),
.sel(s_logisimNet157));
BitSelector
#(.nrOfExtendedBits(65),
.nrOfInputBits(64),
.nrOfselBits(6))
PLEXERS_62
(.dataIn(s_logisimBus187[63:0]),
.dataOut(s_logisimNet107),
.sel(s_logisimBus22[5:0]));
Multiplexer_bus_2
#(.nrOfBits(6))
PLEXERS_63
(.enable(1'b1),
.muxIn_0(s_logisimBus188[5:0]),
.muxIn_1(s_logisimBus47[5:0]),
.muxOut(s_logisimBus16[5:0]),
.sel(s_logisimNet107));
Multiplexer_bus_2
#(.nrOfBits(6))
PLEXERS_64
(.enable(1'b1),
.muxIn_0(s_logisimBus191[5:0]),
.muxIn_1(s_logisimBus161[5:0]),
.muxOut(s_logisimBus144[5:0]),
.sel(s_logisimNet85));
BitSelector
#(.nrOfExtendedBits(65),
.nrOfInputBits(64),
.nrOfselBits(6))
PLEXERS_65
(.dataIn(s_logisimBus187[63:0]),
.dataOut(s_logisimNet15),
.sel(s_logisimBus113[5:0]));
Multiplexer_bus_2
#(.nrOfBits(6))
PLEXERS_66
(.enable(1'b1),
.muxIn_0(s_logisimBus16[5:0]),
.muxIn_1(s_logisimBus140[5:0]),
.muxOut(s_logisimBus95[5:0]),
.sel(s_logisimNet15));
BitSelector
#(.nrOfExtendedBits(65),
.nrOfInputBits(64),
.nrOfselBits(6))
PLEXERS_67
(.dataIn(s_logisimBus187[63:0]),
.dataOut(s_logisimNet61),
.sel(s_logisimBus160[5:0]));
Multiplexer_bus_2
#(.nrOfBits(6))
PLEXERS_68
(.enable(1'b1),
.muxIn_0(s_logisimBus95[5:0]),
.muxIn_1(s_logisimBus184[5:0]),
.muxOut(s_logisimBus53[5:0]),
.sel(s_logisimNet61));
BitSelector
#(.nrOfExtendedBits(65),
.nrOfInputBits(64),
.nrOfselBits(6))
PLEXERS_69
(.dataIn(s_logisimBus187[63:0]),
.dataOut(s_logisimNet180),
.sel(s_logisimBus92[5:0]));
Multiplexer_bus_2
#(.nrOfBits(6))
PLEXERS_70
(.enable(1'b1),
.muxIn_0(s_logisimBus53[5:0]),
.muxIn_1(s_logisimBus21[5:0]),
.muxOut(s_logisimBus77[5:0]),
.sel(s_logisimNet180));
BitSelector
#(.nrOfExtendedBits(65),
.nrOfInputBits(64),
.nrOfselBits(6))
PLEXERS_71
(.dataIn(s_logisimBus187[63:0]),
.dataOut(s_logisimNet14),
.sel(s_logisimBus111[5:0]));
Multiplexer_bus_2
#(.nrOfBits(6))
PLEXERS_72
(.enable(1'b1),
.muxIn_0(s_logisimBus77[5:0]),
.muxIn_1(s_logisimBus137[5:0]),
.muxOut(s_logisimBus75[5:0]),
.sel(s_logisimNet14));
BitSelector
#(.nrOfExtendedBits(65),
.nrOfInputBits(64),
.nrOfselBits(6))
PLEXERS_73
(.dataIn(s_logisimBus187[63:0]),
.dataOut(s_logisimNet154),
.sel(s_logisimBus65[5:0]));
Multiplexer_bus_2
#(.nrOfBits(6))
PLEXERS_74
(.enable(1'b1),
.muxIn_0(s_logisimBus75[5:0]),
.muxIn_1(s_logisimBus90[5:0]),
.muxOut(s_logisimBus189[5:0]),
.sel(s_logisimNet154));
BitSelector
#(.nrOfExtendedBits(65),
.nrOfInputBits(64),
.nrOfselBits(6))
PLEXERS_75
(.dataIn(s_logisimBus187[63:0]),
.dataOut(s_logisimNet37),
.sel(s_logisimBus134[5:0]));
Multiplexer_bus_2
#(.nrOfBits(6))
PLEXERS_76
(.enable(1'b1),
.muxIn_0(s_logisimBus189[5:0]),
.muxIn_1(s_logisimBus68[5:0]),
.muxOut(s_logisimBus100[5:0]),
.sel(s_logisimNet37));
BitSelector
#(.nrOfExtendedBits(65),
.nrOfInputBits(64),
.nrOfselBits(6))
PLEXERS_77
(.dataIn(s_logisimBus187[63:0]),
.dataOut(s_logisimNet176),
.sel(s_logisimBus86[5:0]));
Multiplexer_bus_2
#(.nrOfBits(6))
PLEXERS_78
(.enable(1'b1),
.muxIn_0(s_logisimBus100[5:0]),
.muxIn_1(s_logisimBus17[5:0]),
.muxOut(s_logisimBus156[5:0]),
.sel(s_logisimNet176));
BitSelector
#(.nrOfExtendedBits(65),
.nrOfInputBits(64),
.nrOfselBits(6))
PLEXERS_79
(.dataIn(s_logisimBus187[63:0]),
.dataOut(s_logisimNet38),
.sel(s_logisimBus138[5:0]));
BitSelector
#(.nrOfExtendedBits(65),
.nrOfInputBits(64),
.nrOfselBits(6))
PLEXERS_80
(.dataIn(s_logisimBus187[63:0]),
.dataOut(s_logisimNet105),
.sel(s_logisimBus19[5:0]));
Multiplexer_bus_2
#(.nrOfBits(6))
PLEXERS_81
(.enable(1'b1),
.muxIn_0(s_logisimBus156[5:0]),
.muxIn_1(s_logisimBus42[5:0]),
.muxOut(s_logisimBus11[5:0]),
.sel(s_logisimNet105));
BitSelector
#(.nrOfExtendedBits(65),
.nrOfInputBits(64),
.nrOfselBits(6))
PLEXERS_82
(.dataIn(s_logisimBus187[63:0]),
.dataOut(s_logisimNet5),
.sel(s_logisimBus120[5:0]));
Multiplexer_bus_2
#(.nrOfBits(6))
PLEXERS_83
(.enable(1'b1),
.muxIn_0(s_logisimBus11[5:0]),
.muxIn_1(s_logisimBus147[5:0]),
.muxOut(s_logisimBus51[5:0]),
.sel(s_logisimNet5));
Multiplexer_bus_2
#(.nrOfBits(6))
PLEXERS_84
(.enable(1'b1),
.muxIn_0(s_logisimBus144[5:0]),
.muxIn_1(s_logisimBus112[5:0]),
.muxOut(s_logisimBus97[5:0]),
.sel(s_logisimNet38));
BitSelector
#(.nrOfExtendedBits(65),
.nrOfInputBits(64),
.nrOfselBits(6))
PLEXERS_85
(.dataIn(s_logisimBus187[63:0]),
.dataOut(s_logisimNet81),
.sel(s_logisimBus194[5:0]));
Multiplexer_bus_2
#(.nrOfBits(6))
PLEXERS_86
(.enable(1'b1),
.muxIn_0(s_logisimBus51[5:0]),
.muxIn_1(s_logisimBus123[5:0]),
.muxOut(s_logisimBus72[5:0]),
.sel(s_logisimNet81));
BitSelector
#(.nrOfExtendedBits(65),
.nrOfInputBits(64),
.nrOfselBits(6))
PLEXERS_87
(.dataIn(s_logisimBus187[63:0]),
.dataOut(s_logisimNet32),
.sel(s_logisimBus145[5:0]));
Multiplexer_bus_2
#(.nrOfBits(8))
PLEXERS_88
(.enable(1'b1),
.muxIn_0(s_logisimBus72[7:0]),
.muxIn_1(s_logisimBus76[7:0]),
.muxOut(s_logisimBus8[7:0]),
.sel(s_logisimNet32));
BitSelector
#(.nrOfExtendedBits(65),
.nrOfInputBits(64),
.nrOfselBits(6))
PLEXERS_89
(.dataIn(s_logisimBus187[63:0]),
.dataOut(s_logisimNet179),
.sel(s_logisimBus91[5:0]));
Multiplexer_bus_2
#(.nrOfBits(6))
PLEXERS_90
(.enable(1'b1),
.muxIn_0(s_logisimBus97[5:0]),
.muxIn_1(s_logisimBus67[5:0]),
.muxOut(s_logisimBus114[5:0]),
.sel(s_logisimNet179));
BitSelector
#(.nrOfExtendedBits(65),
.nrOfInputBits(64),
.nrOfselBits(6))
PLEXERS_91
(.dataIn(s_logisimBus187[63:0]),
.dataOut(s_logisimNet59),
.sel(s_logisimBus159[5:0]));
Multiplexer_bus_2
#(.nrOfBits(6))
PLEXERS_92
(.enable(1'b1),
.muxIn_0(s_logisimBus114[5:0]),
.muxIn_1(s_logisimBus135[5:0]),
.muxOut(s_logisimBus119[5:0]),
.sel(s_logisimNet59));
BitSelector
#(.nrOfExtendedBits(65),
.nrOfInputBits(64),
.nrOfselBits(6))
PLEXERS_93
(.dataIn(s_logisimBus187[63:0]),
.dataOut(s_logisimNet10),
.sel(s_logisimBus108[5:0]));
Multiplexer_bus_2
#(.nrOfBits(6))
PLEXERS_94
(.enable(1'b1),
.muxIn_0(s_logisimBus119[5:0]),
.muxIn_1(s_logisimBus87[5:0]),
.muxOut(s_logisimBus103[5:0]),
.sel(s_logisimNet10));
BitSelector
#(.nrOfExtendedBits(65),
.nrOfInputBits(64),
.nrOfselBits(6))
PLEXERS_95
(.dataIn(s_logisimBus187[63:0]),
.dataOut(s_logisimNet127),
.sel(s_logisimBus41[5:0]));
Multiplexer_bus_2
#(.nrOfBits(6))
PLEXERS_96
(.enable(1'b1),
.muxIn_0(s_logisimBus103[5:0]),
.muxIn_1(s_logisimBus18[5:0]),
.muxOut(s_logisimBus195[5:0]),
.sel(s_logisimNet127));
endmodule