/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
CLOO
**
**
**
*****************************************************************************/
module
CLOO(
a,
res_high,
res_low
);
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
[31:0]
a;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
[31:0]
res_high;
output
[31:0]
res_low;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
[5:0]
s_logisimBus0;
wire
[7:0]
s_logisimBus1;
wire
[5:0]
s_logisimBus12;
wire
[5:0]
s_logisimBus14;
wire
[31:0]
s_logisimBus16;
wire
[5:0]
s_logisimBus19;
wire
[3:0]
s_logisimBus25;
wire
[31:0]
s_logisimBus26;
wire
[5:0]
s_logisimBus27;
wire
[5:0]
s_logisimBus28;
wire
[5:0]
s_logisimBus29;
wire
[5:0]
s_logisimBus3;
wire
[5:0]
s_logisimBus31;
wire
[31:0]
s_logisimBus32;
wire
[15:0]
s_logisimBus33;
wire
[1:0]
s_logisimBus34;
wire
[5:0]
s_logisimBus35;
wire
[5:0]
s_logisimBus36;
wire
[15:0]
s_logisimBus37;
wire
[5:0]
s_logisimBus38;
wire
[7:0]
s_logisimBus39;
wire
[5:0]
s_logisimBus40;
wire
[3:0]
s_logisimBus41;
wire
[5:0]
s_logisimBus42;
wire
[1:0]
s_logisimBus43;
wire
[5:0]
s_logisimBus44;
wire
[5:0]
s_logisimBus5;
wire
[5:0]
s_logisimBus7;
wire
[5:0]
s_logisimBus9;
wire
s_logisimNet10;
wire
s_logisimNet11;
wire
s_logisimNet15;
wire
s_logisimNet17;
wire
s_logisimNet21;
wire
s_logisimNet22;
wire
s_logisimNet23;
wire
s_logisimNet24;
wire
s_logisimNet45;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
all
input
connections
are
defined
**
*******************************************************************************/
assign
s_logisimBus16[31:0]
=
a;
/*******************************************************************************
**
Here
all
output
connections
are
defined
**
*******************************************************************************/
assign
res_high
=
s_logisimBus32[31:0];
assign
res_low
=
s_logisimBus26[31:0];
/*******************************************************************************
**
Here
all
in-lined
components
are
defined
**
*******************************************************************************/
assign
s_logisimBus35[5:0]
=
{2'b00,
4'h0};
assign
s_logisimBus32[31:0]
=
32'h00000000;
assign
s_logisimBus26[0]
=
s_logisimBus29[0];
assign
s_logisimBus26[1]
=
s_logisimBus29[1];
assign
s_logisimBus26[2]
=
s_logisimBus29[2];
assign
s_logisimBus26[3]
=
s_logisimBus29[3];
assign
s_logisimBus26[4]
=
s_logisimBus29[4];
assign
s_logisimBus26[5]
=
s_logisimBus29[5];
assign
s_logisimBus26[6]
=
1'b0;
assign
s_logisimBus26[7]
=
1'b0;
assign
s_logisimBus26[8]
=
1'b0;
assign
s_logisimBus26[9]
=
1'b0;
assign
s_logisimBus26[10]
=
1'b0;
assign
s_logisimBus26[11]
=
1'b0;
assign
s_logisimBus26[12]
=
1'b0;
assign
s_logisimBus26[13]
=
1'b0;
assign
s_logisimBus26[14]
=
1'b0;
assign
s_logisimBus26[15]
=
1'b0;
assign
s_logisimBus26[16]
=
1'b0;
assign
s_logisimBus26[17]
=
1'b0;
assign
s_logisimBus26[18]
=
1'b0;
assign
s_logisimBus26[19]
=
1'b0;
assign
s_logisimBus26[20]
=
1'b0;
assign
s_logisimBus26[21]
=
1'b0;
assign
s_logisimBus26[22]
=
1'b0;
assign
s_logisimBus26[23]
=
1'b0;
assign
s_logisimBus26[24]
=
1'b0;
assign
s_logisimBus26[25]
=
1'b0;
assign
s_logisimBus26[26]
=
1'b0;
assign
s_logisimBus26[27]
=
1'b0;
assign
s_logisimBus26[28]
=
1'b0;
assign
s_logisimBus26[29]
=
1'b0;
assign
s_logisimBus26[30]
=
1'b0;
assign
s_logisimBus26[31]
=
1'b0;
assign
s_logisimBus9[5:0]
=
{2'b00,
4'h0};
assign
s_logisimBus36[5:0]
=
{2'b00,
4'h1};
assign
s_logisimBus37[15:0]
=
16'hFFFF;
assign
s_logisimBus38[5:0]
=
{2'b00,
4'h8};
assign
s_logisimBus39[7:0]
=
8'hFF;
assign
s_logisimBus40[5:0]
=
{2'b00,
4'h4};
assign
s_logisimBus41[3:0]
=
4'hF;
assign
s_logisimBus42[5:0]
=
{2'b00,
4'h2};
assign
s_logisimBus43[1:0]
=
2'b11;
assign
s_logisimBus44[5:0]
=
{2'b00,
4'h1};
assign
s_logisimNet45
=
1'b1;
/*******************************************************************************
**
Here
all
normal
components
are
defined
**
*******************************************************************************/
Multiplexer_bus_2
#(.nrOfBits(16))
PLEXERS_1
(.enable(1'b1),
.muxIn_0(s_logisimBus16[31:16]),
.muxIn_1(s_logisimBus16[15:0]),
.muxOut(s_logisimBus33[15:0]),
.sel(s_logisimNet17));
Multiplexer_bus_2
#(.nrOfBits(6))
PLEXERS_2
(.enable(1'b1),
.muxIn_0(s_logisimBus9[5:0]),
.muxIn_1(s_logisimBus3[5:0]),
.muxOut(s_logisimBus27[5:0]),
.sel(s_logisimNet17));
Multiplexer_bus_2
#(.nrOfBits(8))
PLEXERS_3
(.enable(1'b1),
.muxIn_0(s_logisimBus33[15:8]),
.muxIn_1(s_logisimBus33[7:0]),
.muxOut(s_logisimBus1[7:0]),
.sel(s_logisimNet21));
Multiplexer_bus_2
#(.nrOfBits(6))
PLEXERS_4
(.enable(1'b1),
.muxIn_0(s_logisimBus27[5:0]),
.muxIn_1(s_logisimBus31[5:0]),
.muxOut(s_logisimBus14[5:0]),
.sel(s_logisimNet21));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_5
(.enable(1'b1),
.muxIn_0(s_logisimBus1[7:4]),
.muxIn_1(s_logisimBus1[3:0]),
.muxOut(s_logisimBus25[3:0]),
.sel(s_logisimNet22));
Multiplexer_bus_2
#(.nrOfBits(6))
PLEXERS_6
(.enable(1'b1),
.muxIn_0(s_logisimBus14[5:0]),
.muxIn_1(s_logisimBus28[5:0]),
.muxOut(s_logisimBus0[5:0]),
.sel(s_logisimNet22));
Multiplexer_bus_2
#(.nrOfBits(2))
PLEXERS_7
(.enable(1'b1),
.muxIn_0(s_logisimBus25[3:2]),
.muxIn_1(s_logisimBus25[1:0]),
.muxOut(s_logisimBus34[1:0]),
.sel(s_logisimNet11));
Multiplexer_bus_2
#(.nrOfBits(6))
PLEXERS_8
(.enable(1'b1),
.muxIn_0(s_logisimBus0[5:0]),
.muxIn_1(s_logisimBus19[5:0]),
.muxOut(s_logisimBus12[5:0]),
.sel(s_logisimNet11));
Multiplexer_2
PLEXERS_9
(.enable(1'b1),
.muxIn_0(s_logisimBus34[1]),
.muxIn_1(s_logisimBus34[0]),
.muxOut(s_logisimNet23),
.sel(s_logisimNet10));
Multiplexer_bus_2
#(.nrOfBits(6))
PLEXERS_10
(.enable(1'b1),
.muxIn_0(s_logisimBus12[5:0]),
.muxIn_1(s_logisimBus5[5:0]),
.muxOut(s_logisimBus7[5:0]),
.sel(s_logisimNet10));
Adder
#(.extendedBits(7),
.nrOfBits(6))
ARITH_11
(.carryIn(s_logisimNet23),
.carryOut(),
.dataA(s_logisimBus35[5:0]),
.dataB(s_logisimBus7[5:0]),
.result(s_logisimBus29[5:0]));
Adder
#(.extendedBits(7),
.nrOfBits(6))
ARITH_12
(.carryIn(1'b0),
.carryOut(),
.dataA(s_logisimBus9[5:0]),
.dataB(s_logisimBus36[5:0]),
.result(s_logisimBus3[5:0]));
Comparator
#(.nrOfBits(16),
.twosComplement(0))
ARITH_13
(.aEqualsB(s_logisimNet17),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus16[31:16]),
.dataB(s_logisimBus37[15:0]));
Adder
#(.extendedBits(7),
.nrOfBits(6))
ARITH_14
(.carryIn(1'b0),
.carryOut(),
.dataA(s_logisimBus27[5:0]),
.dataB(s_logisimBus38[5:0]),
.result(s_logisimBus31[5:0]));
Comparator
#(.nrOfBits(8),
.twosComplement(0))
ARITH_15
(.aEqualsB(s_logisimNet21),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus33[15:8]),
.dataB(s_logisimBus39[7:0]));
Adder
#(.extendedBits(7),
.nrOfBits(6))
ARITH_16
(.carryIn(1'b0),
.carryOut(),
.dataA(s_logisimBus14[5:0]),
.dataB(s_logisimBus40[5:0]),
.result(s_logisimBus28[5:0]));
Comparator
#(.nrOfBits(4),
.twosComplement(0))
ARITH_17
(.aEqualsB(s_logisimNet22),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus1[7:4]),
.dataB(s_logisimBus41[3:0]));
Adder
#(.extendedBits(7),
.nrOfBits(6))
ARITH_18
(.carryIn(1'b0),
.carryOut(),
.dataA(s_logisimBus0[5:0]),
.dataB(s_logisimBus42[5:0]),
.result(s_logisimBus19[5:0]));
Comparator
#(.nrOfBits(2),
.twosComplement(0))
ARITH_19
(.aEqualsB(s_logisimNet11),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus25[3:2]),
.dataB(s_logisimBus43[1:0]));
Adder
#(.extendedBits(7),
.nrOfBits(6))
ARITH_20
(.carryIn(1'b0),
.carryOut(),
.dataA(s_logisimBus12[5:0]),
.dataB(s_logisimBus44[5:0]),
.result(s_logisimBus5[5:0]));
BitComparator
#(.twosComplement(0))
ARITH_21
(.aEqualsB(s_logisimNet10),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus34[1]),
.dataB(s_logisimNet45));
endmodule