/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
main
**
**
**
*****************************************************************************/
module
main(
InstDone,
Jen,
Jin,
Jout,
PC,
R1,
R10,
R11,
R12,
R13,
R14,
R15,
R16,
R17,
R18,
R19,
R2,
R20,
R21,
R22,
R23,
R24,
R25,
R26,
R27,
R28,
R29,
R3,
R30,
R31,
R4,
R5,
R6,
R7,
R8,
R9,
clk,
rst
);
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
Jen;
input
[31:0]
Jin;
input
clk;
input
rst;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
InstDone;
output
[31:0]
Jout;
output
[8:0]
PC;
output
[31:0]
R1;
output
[31:0]
R10;
output
[31:0]
R11;
output
[31:0]
R12;
output
[31:0]
R13;
output
[31:0]
R14;
output
[31:0]
R15;
output
[31:0]
R16;
output
[31:0]
R17;
output
[31:0]
R18;
output
[31:0]
R19;
output
[31:0]
R2;
output
[31:0]
R20;
output
[31:0]
R21;
output
[31:0]
R22;
output
[31:0]
R23;
output
[31:0]
R24;
output
[31:0]
R25;
output
[31:0]
R26;
output
[31:0]
R27;
output
[31:0]
R28;
output
[31:0]
R29;
output
[31:0]
R3;
output
[31:0]
R30;
output
[31:0]
R31;
output
[31:0]
R4;
output
[31:0]
R5;
output
[31:0]
R6;
output
[31:0]
R7;
output
[31:0]
R8;
output
[31:0]
R9;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
[4:0]
s_logisimBus0;
wire
[31:0]
s_logisimBus1;
wire
[8:0]
s_logisimBus10;
wire
[31:0]
s_logisimBus100;
wire
[31:0]
s_logisimBus101;
wire
[31:0]
s_logisimBus102;
wire
[31:0]
s_logisimBus103;
wire
[31:0]
s_logisimBus104;
wire
[31:0]
s_logisimBus105;
wire
[31:0]
s_logisimBus106;
wire
[31:0]
s_logisimBus107;
wire
[31:0]
s_logisimBus108;
wire
[31:0]
s_logisimBus109;
wire
[31:0]
s_logisimBus110;
wire
[3:0]
s_logisimBus112;
wire
[31:0]
s_logisimBus13;
wire
[31:0]
s_logisimBus15;
wire
[8:0]
s_logisimBus16;
wire
[4:0]
s_logisimBus18;
wire
[31:0]
s_logisimBus2;
wire
[4:0]
s_logisimBus20;
wire
[31:0]
s_logisimBus21;
wire
[5:0]
s_logisimBus22;
wire
[4:0]
s_logisimBus24;
wire
[31:0]
s_logisimBus27;
wire
[31:0]
s_logisimBus28;
wire
[31:0]
s_logisimBus29;
wire
[4:0]
s_logisimBus3;
wire
[31:0]
s_logisimBus30;
wire
[8:0]
s_logisimBus31;
wire
[4:0]
s_logisimBus32;
wire
[8:0]
s_logisimBus33;
wire
[8:0]
s_logisimBus34;
wire
[31:0]
s_logisimBus35;
wire
[31:0]
s_logisimBus36;
wire
[8:0]
s_logisimBus38;
wire
[4:0]
s_logisimBus4;
wire
[8:0]
s_logisimBus40;
wire
[31:0]
s_logisimBus41;
wire
[4:0]
s_logisimBus42;
wire
[8:0]
s_logisimBus44;
wire
[8:0]
s_logisimBus46;
wire
[31:0]
s_logisimBus47;
wire
[31:0]
s_logisimBus48;
wire
[31:0]
s_logisimBus49;
wire
[4:0]
s_logisimBus5;
wire
[4:0]
s_logisimBus51;
wire
[8:0]
s_logisimBus52;
wire
[31:0]
s_logisimBus53;
wire
[4:0]
s_logisimBus56;
wire
[5:0]
s_logisimBus58;
wire
[31:0]
s_logisimBus59;
wire
[15:0]
s_logisimBus6;
wire
[31:0]
s_logisimBus61;
wire
[31:0]
s_logisimBus62;
wire
[31:0]
s_logisimBus63;
wire
[31:0]
s_logisimBus65;
wire
[4:0]
s_logisimBus66;
wire
[31:0]
s_logisimBus68;
wire
[31:0]
s_logisimBus69;
wire
[4:0]
s_logisimBus7;
wire
[31:0]
s_logisimBus71;
wire
[31:0]
s_logisimBus72;
wire
[8:0]
s_logisimBus76;
wire
[31:0]
s_logisimBus79;
wire
[4:0]
s_logisimBus8;
wire
[31:0]
s_logisimBus80;
wire
[31:0]
s_logisimBus81;
wire
[31:0]
s_logisimBus82;
wire
[31:0]
s_logisimBus83;
wire
[31:0]
s_logisimBus84;
wire
[31:0]
s_logisimBus85;
wire
[31:0]
s_logisimBus86;
wire
[31:0]
s_logisimBus87;
wire
[31:0]
s_logisimBus88;
wire
[31:0]
s_logisimBus89;
wire
[4:0]
s_logisimBus9;
wire
[31:0]
s_logisimBus90;
wire
[31:0]
s_logisimBus91;
wire
[31:0]
s_logisimBus92;
wire
[31:0]
s_logisimBus93;
wire
[31:0]
s_logisimBus94;
wire
[31:0]
s_logisimBus95;
wire
[31:0]
s_logisimBus96;
wire
[31:0]
s_logisimBus97;
wire
[31:0]
s_logisimBus98;
wire
[31:0]
s_logisimBus99;
wire
s_logisimNet11;
wire
s_logisimNet111;
wire
s_logisimNet12;
wire
s_logisimNet14;
wire
s_logisimNet17;
wire
s_logisimNet19;
wire
s_logisimNet23;
wire
s_logisimNet25;
wire
s_logisimNet26;
wire
s_logisimNet37;
wire
s_logisimNet39;
wire
s_logisimNet43;
wire
s_logisimNet45;
wire
s_logisimNet50;
wire
s_logisimNet54;
wire
s_logisimNet55;
wire
s_logisimNet57;
wire
s_logisimNet60;
wire
s_logisimNet64;
wire
s_logisimNet67;
wire
s_logisimNet70;
wire
s_logisimNet77;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
all
input
connections
are
defined
**
*******************************************************************************/
assign
s_logisimBus69[31:0]
=
Jin;
assign
s_logisimNet11
=
Jen;
assign
s_logisimNet111
=
clk;
assign
s_logisimNet77
=
rst;
/*******************************************************************************
**
Here
all
output
connections
are
defined
**
*******************************************************************************/
assign
InstDone
=
s_logisimNet12;
assign
Jout
=
s_logisimBus79[31:0];
assign
PC
=
s_logisimBus10[8:0];
assign
R1
=
s_logisimBus80[31:0];
assign
R10
=
s_logisimBus89[31:0];
assign
R11
=
s_logisimBus90[31:0];
assign
R12
=
s_logisimBus91[31:0];
assign
R13
=
s_logisimBus92[31:0];
assign
R14
=
s_logisimBus93[31:0];
assign
R15
=
s_logisimBus94[31:0];
assign
R16
=
s_logisimBus95[31:0];
assign
R17
=
s_logisimBus96[31:0];
assign
R18
=
s_logisimBus97[31:0];
assign
R19
=
s_logisimBus98[31:0];
assign
R2
=
s_logisimBus81[31:0];
assign
R20
=
s_logisimBus99[31:0];
assign
R21
=
s_logisimBus100[31:0];
assign
R22
=
s_logisimBus101[31:0];
assign
R23
=
s_logisimBus102[31:0];
assign
R24
=
s_logisimBus103[31:0];
assign
R25
=
s_logisimBus104[31:0];
assign
R26
=
s_logisimBus105[31:0];
assign
R27
=
s_logisimBus106[31:0];
assign
R28
=
s_logisimBus107[31:0];
assign
R29
=
s_logisimBus108[31:0];
assign
R3
=
s_logisimBus82[31:0];
assign
R30
=
s_logisimBus109[31:0];
assign
R31
=
s_logisimBus110[31:0];
assign
R4
=
s_logisimBus83[31:0];
assign
R5
=
s_logisimBus84[31:0];
assign
R6
=
s_logisimBus85[31:0];
assign
R7
=
s_logisimBus86[31:0];
assign
R8
=
s_logisimBus87[31:0];
assign
R9
=
s_logisimBus88[31:0];
/*******************************************************************************
**
Here
all
in-lined
components
are
defined
**
*******************************************************************************/
assign
s_logisimBus46[8:0]
=
{1'b0,
8'h01};
assign
s_logisimBus47[0]
=
s_logisimBus6[0];
assign
s_logisimBus47[1]
=
s_logisimBus6[1];
assign
s_logisimBus47[2]
=
s_logisimBus6[2];
assign
s_logisimBus47[3]
=
s_logisimBus6[3];
assign
s_logisimBus47[4]
=
s_logisimBus6[4];
assign
s_logisimBus47[5]
=
s_logisimBus6[5];
assign
s_logisimBus47[6]
=
s_logisimBus6[6];
assign
s_logisimBus47[7]
=
s_logisimBus6[7];
assign
s_logisimBus47[8]
=
s_logisimBus6[8];
assign
s_logisimBus47[9]
=
s_logisimBus6[9];
assign
s_logisimBus47[10]
=
s_logisimBus6[10];
assign
s_logisimBus47[11]
=
s_logisimBus6[11];
assign
s_logisimBus47[12]
=
s_logisimBus6[12];
assign
s_logisimBus47[13]
=
s_logisimBus6[13];
assign
s_logisimBus47[14]
=
s_logisimBus6[14];
assign
s_logisimBus47[15]
=
s_logisimBus6[15];
assign
s_logisimBus47[16]
=
s_logisimBus6[15];
assign
s_logisimBus47[17]
=
s_logisimBus6[15];
assign
s_logisimBus47[18]
=
s_logisimBus6[15];
assign
s_logisimBus47[19]
=
s_logisimBus6[15];
assign
s_logisimBus47[20]
=
s_logisimBus6[15];
assign
s_logisimBus47[21]
=
s_logisimBus6[15];
assign
s_logisimBus47[22]
=
s_logisimBus6[15];
assign
s_logisimBus47[23]
=
s_logisimBus6[15];
assign
s_logisimBus47[24]
=
s_logisimBus6[15];
assign
s_logisimBus47[25]
=
s_logisimBus6[15];
assign
s_logisimBus47[26]
=
s_logisimBus6[15];
assign
s_logisimBus47[27]
=
s_logisimBus6[15];
assign
s_logisimBus47[28]
=
s_logisimBus6[15];
assign
s_logisimBus47[29]
=
s_logisimBus6[15];
assign
s_logisimBus47[30]
=
s_logisimBus6[15];
assign
s_logisimBus47[31]
=
s_logisimBus6[15];
assign
s_logisimBus35[0]
=
s_logisimBus32[0];
assign
s_logisimBus35[1]
=
s_logisimBus32[1];
assign
s_logisimBus35[2]
=
s_logisimBus32[2];
assign
s_logisimBus35[3]
=
s_logisimBus32[3];
assign
s_logisimBus35[4]
=
s_logisimBus32[4];
assign
s_logisimBus35[5]
=
1'b0;
assign
s_logisimBus35[6]
=
1'b0;
assign
s_logisimBus35[7]
=
1'b0;
assign
s_logisimBus35[8]
=
1'b0;
assign
s_logisimBus35[9]
=
1'b0;
assign
s_logisimBus35[10]
=
1'b0;
assign
s_logisimBus35[11]
=
1'b0;
assign
s_logisimBus35[12]
=
1'b0;
assign
s_logisimBus35[13]
=
1'b0;
assign
s_logisimBus35[14]
=
1'b0;
assign
s_logisimBus35[15]
=
1'b0;
assign
s_logisimBus35[16]
=
1'b0;
assign
s_logisimBus35[17]
=
1'b0;
assign
s_logisimBus35[18]
=
1'b0;
assign
s_logisimBus35[19]
=
1'b0;
assign
s_logisimBus35[20]
=
1'b0;
assign
s_logisimBus35[21]
=
1'b0;
assign
s_logisimBus35[22]
=
1'b0;
assign
s_logisimBus35[23]
=
1'b0;
assign
s_logisimBus35[24]
=
1'b0;
assign
s_logisimBus35[25]
=
1'b0;
assign
s_logisimBus35[26]
=
1'b0;
assign
s_logisimBus35[27]
=
1'b0;
assign
s_logisimBus35[28]
=
1'b0;
assign
s_logisimBus35[29]
=
1'b0;
assign
s_logisimBus35[30]
=
1'b0;
assign
s_logisimBus35[31]
=
1'b0;
assign
s_logisimBus29[0]
=
s_logisimBus52[0];
assign
s_logisimBus29[1]
=
s_logisimBus52[1];
assign
s_logisimBus29[2]
=
s_logisimBus52[2];
assign
s_logisimBus29[3]
=
s_logisimBus52[3];
assign
s_logisimBus29[4]
=
s_logisimBus52[4];
assign
s_logisimBus29[5]
=
s_logisimBus52[5];
assign
s_logisimBus29[6]
=
s_logisimBus52[6];
assign
s_logisimBus29[7]
=
s_logisimBus52[7];
assign
s_logisimBus29[8]
=
s_logisimBus52[8];
assign
s_logisimBus29[9]
=
s_logisimBus52[8];
assign
s_logisimBus29[10]
=
s_logisimBus52[8];
assign
s_logisimBus29[11]
=
s_logisimBus52[8];
assign
s_logisimBus29[12]
=
s_logisimBus52[8];
assign
s_logisimBus29[13]
=
s_logisimBus52[8];
assign
s_logisimBus29[14]
=
s_logisimBus52[8];
assign
s_logisimBus29[15]
=
s_logisimBus52[8];
assign
s_logisimBus29[16]
=
s_logisimBus52[8];
assign
s_logisimBus29[17]
=
s_logisimBus52[8];
assign
s_logisimBus29[18]
=
s_logisimBus52[8];
assign
s_logisimBus29[19]
=
s_logisimBus52[8];
assign
s_logisimBus29[20]
=
s_logisimBus52[8];
assign
s_logisimBus29[21]
=
s_logisimBus52[8];
assign
s_logisimBus29[22]
=
s_logisimBus52[8];
assign
s_logisimBus29[23]
=
s_logisimBus52[8];
assign
s_logisimBus29[24]
=
s_logisimBus52[8];
assign
s_logisimBus29[25]
=
s_logisimBus52[8];
assign
s_logisimBus29[26]
=
s_logisimBus52[8];
assign
s_logisimBus29[27]
=
s_logisimBus52[8];
assign
s_logisimBus29[28]
=
s_logisimBus52[8];
assign
s_logisimBus29[29]
=
s_logisimBus52[8];
assign
s_logisimBus29[30]
=
s_logisimBus52[8];
assign
s_logisimBus29[31]
=
s_logisimBus52[8];
assign
s_logisimBus51[4:0]
=
{1'b0,
4'h0};
assign
s_logisimBus28[0]
=
s_logisimBus5[0];
assign
s_logisimBus28[1]
=
s_logisimBus5[1];
assign
s_logisimBus28[2]
=
s_logisimBus5[2];
assign
s_logisimBus28[3]
=
s_logisimBus5[3];
assign
s_logisimBus28[4]
=
s_logisimBus5[4];
assign
s_logisimBus28[5]
=
1'b0;
assign
s_logisimBus28[6]
=
1'b0;
assign
s_logisimBus28[7]
=
1'b0;
assign
s_logisimBus28[8]
=
1'b0;
assign
s_logisimBus28[9]
=
1'b0;
assign
s_logisimBus28[10]
=
1'b0;
assign
s_logisimBus28[11]
=
1'b0;
assign
s_logisimBus28[12]
=
1'b0;
assign
s_logisimBus28[13]
=
1'b0;
assign
s_logisimBus28[14]
=
1'b0;
assign
s_logisimBus28[15]
=
1'b0;
assign
s_logisimBus28[16]
=
1'b0;
assign
s_logisimBus28[17]
=
1'b0;
assign
s_logisimBus28[18]
=
1'b0;
assign
s_logisimBus28[19]
=
1'b0;
assign
s_logisimBus28[20]
=
1'b0;
assign
s_logisimBus28[21]
=
1'b0;
assign
s_logisimBus28[22]
=
1'b0;
assign
s_logisimBus28[23]
=
1'b0;
assign
s_logisimBus28[24]
=
1'b0;
assign
s_logisimBus28[25]
=
1'b0;
assign
s_logisimBus28[26]
=
1'b0;
assign
s_logisimBus28[27]
=
1'b0;
assign
s_logisimBus28[28]
=
1'b0;
assign
s_logisimBus28[29]
=
1'b0;
assign
s_logisimBus28[30]
=
1'b0;
assign
s_logisimBus28[31]
=
1'b0;
assign
s_logisimBus56[4:0]
=
{1'b1,
4'hF};
/*******************************************************************************
**
Here
all
normal
components
are
defined
**
*******************************************************************************/
AND_GATE
#(.BubblesMask(2'b01))
GATES_1
(.input1(s_logisimNet43),
.input2(s_logisimNet70),
.result(s_logisimNet23));
OR_GATE
#(.BubblesMask(2'b00))
GATES_2
(.input1(s_logisimNet23),
.input2(s_logisimNet54),
.result(s_logisimNet17));
AND_GATE
#(.BubblesMask(2'b00))
GATES_3
(.input1(s_logisimNet43),
.input2(s_logisimNet14),
.result(s_logisimNet54));
OR_GATE
#(.BubblesMask(2'b00))
GATES_4
(.input1(s_logisimNet50),
.input2(s_logisimNet55),
.result(s_logisimNet39));
Multiplexer_bus_2
#(.nrOfBits(5))
PLEXERS_5
(.enable(1'b1),
.muxIn_0(s_logisimBus7[4:0]),
.muxIn_1(s_logisimBus24[4:0]),
.muxOut(s_logisimBus3[4:0]),
.sel(s_logisimNet45));
Multiplexer_bus_2
#(.nrOfBits(5))
PLEXERS_6
(.enable(1'b1),
.muxIn_0(s_logisimBus3[4:0]),
.muxIn_1(s_logisimBus42[4:0]),
.muxOut(s_logisimBus8[4:0]),
.sel(s_logisimNet37));
Multiplexer_bus_2
#(.nrOfBits(32))
PLEXERS_7
(.enable(1'b1),
.muxIn_0(s_logisimBus49[31:0]),
.muxIn_1(s_logisimBus59[31:0]),
.muxOut(s_logisimBus1[31:0]),
.sel(s_logisimNet64));
Multiplexer_bus_2
#(.nrOfBits(32))
PLEXERS_8
(.enable(1'b1),
.muxIn_0(s_logisimBus1[31:0]),
.muxIn_1(s_logisimBus29[31:0]),
.muxOut(s_logisimBus63[31:0]),
.sel(s_logisimNet67));
Multiplexer_bus_2
#(.nrOfBits(5))
PLEXERS_9
(.enable(1'b1),
.muxIn_0(s_logisimBus51[4:0]),
.muxIn_1(s_logisimBus66[4:0]),
.muxOut(s_logisimBus0[4:0]),
.sel(s_logisimNet60));
Multiplexer_bus_2
#(.nrOfBits(5))
PLEXERS_10
(.enable(1'b1),
.muxIn_0(s_logisimBus0[4:0]),
.muxIn_1(s_logisimBus56[4:0]),
.muxOut(s_logisimBus5[4:0]),
.sel(s_logisimNet67));
Multiplexer_bus_2
#(.nrOfBits(32))
PLEXERS_11
(.enable(1'b1),
.muxIn_0(s_logisimBus65[31:0]),
.muxIn_1(s_logisimBus68[31:0]),
.muxOut(s_logisimBus27[31:0]),
.sel(s_logisimNet19));
Multiplexer_bus_2
#(.nrOfBits(32))
PLEXERS_12
(.enable(1'b1),
.muxIn_0(s_logisimBus27[31:0]),
.muxIn_1(s_logisimBus48[31:0]),
.muxOut(s_logisimBus61[31:0]),
.sel(s_logisimNet26));
Multiplexer_bus_2
#(.nrOfBits(32))
PLEXERS_13
(.enable(1'b1),
.muxIn_0(s_logisimBus71[31:0]),
.muxIn_1(s_logisimBus65[31:0]),
.muxOut(s_logisimBus21[31:0]),
.sel(s_logisimNet26));
Multiplexer_bus_2
#(.nrOfBits(9))
PLEXERS_14
(.enable(1'b1),
.muxIn_0(s_logisimBus38[8:0]),
.muxIn_1(s_logisimBus44[8:0]),
.muxOut(s_logisimBus34[8:0]),
.sel(s_logisimNet17));
Multiplexer_bus_2
#(.nrOfBits(9))
PLEXERS_15
(.enable(1'b1),
.muxIn_0(s_logisimBus34[8:0]),
.muxIn_1(s_logisimBus68[8:0]),
.muxOut(s_logisimBus31[8:0]),
.sel(s_logisimNet39));
Multiplexer_bus_2
#(.nrOfBits(9))
PLEXERS_16
(.enable(1'b1),
.muxIn_0(s_logisimBus31[8:0]),
.muxIn_1(s_logisimBus71[8:0]),
.muxOut(s_logisimBus33[8:0]),
.sel(s_logisimNet57));
Adder
#(.extendedBits(10),
.nrOfBits(9))
ARITH_17
(.carryIn(1'b0),
.carryOut(),
.dataA(s_logisimBus76[8:0]),
.dataB(s_logisimBus46[8:0]),
.result(s_logisimBus38[8:0]));
Adder
#(.extendedBits(10),
.nrOfBits(9))
ARITH_18
(.carryIn(1'b0),
.carryOut(),
.dataA(s_logisimBus52[8:0]),
.dataB(s_logisimBus68[8:0]),
.result(s_logisimBus44[8:0]));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(9))
MEMORY_19
(.clock(s_logisimNet111),
.clockEnable(1'b1),
.d(s_logisimBus76[8:0]),
.q(s_logisimBus16[8:0]),
.reset(s_logisimNet77),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(32))
MemoryDataReg
(.clock(s_logisimNet111),
.clockEnable(1'b1),
.d(s_logisimBus30[31:0]),
.q(s_logisimBus59[31:0]),
.reset(s_logisimNet77),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(32))
InstructionReg
(.clock(s_logisimNet111),
.clockEnable(1'b1),
.d(s_logisimBus13[31:0]),
.q(s_logisimBus41[31:0]),
.reset(s_logisimNet77),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(5))
MEMORY_22
(.clock(s_logisimNet111),
.clockEnable(1'b1),
.d(s_logisimBus4[4:0]),
.q(s_logisimBus42[4:0]),
.reset(s_logisimNet77),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(5))
MEMORY_23
(.clock(s_logisimNet111),
.clockEnable(1'b1),
.d(s_logisimBus18[4:0]),
.q(s_logisimBus7[4:0]),
.reset(s_logisimNet77),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(5))
MEMORY_24
(.clock(s_logisimNet111),
.clockEnable(1'b1),
.d(s_logisimBus20[4:0]),
.q(s_logisimBus24[4:0]),
.reset(s_logisimNet77),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(32))
MEMORY_25
(.clock(s_logisimNet111),
.clockEnable(1'b1),
.d(s_logisimBus47[31:0]),
.q(s_logisimBus68[31:0]),
.reset(s_logisimNet77),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(32))
MEMORY_26
(.clock(s_logisimNet111),
.clockEnable(1'b1),
.d(s_logisimBus35[31:0]),
.q(s_logisimBus48[31:0]),
.reset(s_logisimNet77),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(5))
MEMORY_27
(.clock(s_logisimNet111),
.clockEnable(1'b1),
.d(s_logisimBus8[4:0]),
.q(s_logisimBus9[4:0]),
.reset(s_logisimNet77),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(5))
MEMORY_28
(.clock(s_logisimNet111),
.clockEnable(1'b1),
.d(s_logisimBus9[4:0]),
.q(s_logisimBus66[4:0]),
.reset(s_logisimNet77),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(9))
MEMORY_29
(.clock(s_logisimNet111),
.clockEnable(1'b1),
.d(s_logisimBus16[8:0]),
.q(s_logisimBus40[8:0]),
.reset(s_logisimNet77),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(32))
A
(.clock(s_logisimNet111),
.clockEnable(1'b1),
.d(s_logisimBus2[31:0]),
.q(s_logisimBus71[31:0]),
.reset(s_logisimNet77),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(32))
B
(.clock(s_logisimNet111),
.clockEnable(1'b1),
.d(s_logisimBus15[31:0]),
.q(s_logisimBus65[31:0]),
.reset(s_logisimNet77),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(32))
MEMORY_32
(.clock(s_logisimNet111),
.clockEnable(1'b1),
.d(s_logisimBus65[31:0]),
.q(s_logisimBus62[31:0]),
.reset(s_logisimNet77),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(9))
MEMORY_33
(.clock(s_logisimNet111),
.clockEnable(1'b1),
.d(s_logisimBus40[8:0]),
.q(s_logisimBus52[8:0]),
.reset(s_logisimNet77),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(32))
MEMORY_34
(.clock(s_logisimNet111),
.clockEnable(1'b1),
.d(s_logisimBus53[31:0]),
.q(s_logisimBus72[31:0]),
.reset(s_logisimNet77),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(32))
MEMORY_35
(.clock(s_logisimNet111),
.clockEnable(1'b1),
.d(s_logisimBus72[31:0]),
.q(s_logisimBus49[31:0]),
.reset(s_logisimNet77),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(9))
MEMORY_36
(.clock(s_logisimNet111),
.clockEnable(1'b1),
.d(s_logisimBus52[8:0]),
.q(s_logisimBus10[8:0]),
.reset(s_logisimNet77),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(9))
pcc
(.clock(s_logisimNet111),
.clockEnable(1'b1),
.d(s_logisimBus33[8:0]),
.q(s_logisimBus76[8:0]),
.reset(s_logisimNet77),
.tick(1'b1));
/*******************************************************************************
**
Here
all
sub-circuits
are
defined
**
*******************************************************************************/
jtag_ram512
Dmem
(.Addr(s_logisimBus72[8:0]),
.Din(s_logisimBus62[31:0]),
.Dout(s_logisimBus30[31:0]),
.Jen(s_logisimNet11),
.Jin(s_logisimBus36[31:0]),
.Jout(s_logisimBus79[31:0]),
.Wen(s_logisimNet25),
.clk(s_logisimNet111));
jtag_ram512
Imem
(.Addr(s_logisimBus76[8:0]),
.Din(32'd0),
.Dout(s_logisimBus13[31:0]),
.Jen(s_logisimNet11),
.Jin(s_logisimBus69[31:0]),
.Jout(s_logisimBus36[31:0]),
.Wen(1'b0),
.clk(s_logisimNet111));
InstructionDecode
x1
(.Instruction(s_logisimBus41[31:0]),
.func(s_logisimBus58[5:0]),
.imm(s_logisimBus6[15:0]),
.opCode(s_logisimBus22[5:0]),
.rd(s_logisimBus20[4:0]),
.rs(s_logisimBus4[4:0]),
.rt(s_logisimBus18[4:0]),
.shmt(s_logisimBus32[4:0]));
regfile
x4
(.Aread0(s_logisimBus18[4:0]),
.Aread1(s_logisimBus4[4:0]),
.Awrite(s_logisimBus5[4:0]),
.Dread0(s_logisimBus2[31:0]),
.Dread1(s_logisimBus15[31:0]),
.Dwrite(s_logisimBus63[31:0]),
.R1(s_logisimBus80[31:0]),
.R10(s_logisimBus89[31:0]),
.R11(s_logisimBus90[31:0]),
.R12(s_logisimBus91[31:0]),
.R13(s_logisimBus92[31:0]),
.R14(s_logisimBus93[31:0]),
.R15(s_logisimBus94[31:0]),
.R16(s_logisimBus95[31:0]),
.R17(s_logisimBus96[31:0]),
.R18(s_logisimBus97[31:0]),
.R19(s_logisimBus98[31:0]),
.R2(s_logisimBus81[31:0]),
.R20(s_logisimBus99[31:0]),
.R21(s_logisimBus100[31:0]),
.R22(s_logisimBus101[31:0]),
.R23(s_logisimBus102[31:0]),
.R24(s_logisimBus103[31:0]),
.R25(s_logisimBus104[31:0]),
.R26(s_logisimBus105[31:0]),
.R27(s_logisimBus106[31:0]),
.R28(s_logisimBus107[31:0]),
.R29(s_logisimBus108[31:0]),
.R3(s_logisimBus82[31:0]),
.R30(s_logisimBus109[31:0]),
.R31(s_logisimBus110[31:0]),
.R4(s_logisimBus83[31:0]),
.R5(s_logisimBus84[31:0]),
.R6(s_logisimBus85[31:0]),
.R7(s_logisimBus86[31:0]),
.R8(s_logisimBus87[31:0]),
.R9(s_logisimBus88[31:0]),
.clk(s_logisimNet111),
.rst(s_logisimNet77));
ALU
x3
(.InstDone(s_logisimNet12),
.a(s_logisimBus21[31:0]),
.aluop(s_logisimBus112[3:0]),
.b(s_logisimBus61[31:0]),
.clk(s_logisimNet111),
.res_high(),
.res_low(s_logisimBus53[31:0]),
.zero(s_logisimNet43));
ControlUnit
ControlUnit_1
(.ALUop(s_logisimBus112[3:0]),
.ALUsrc(s_logisimNet19),
.addi_lw(s_logisimNet37),
.beq(s_logisimNet14),
.branchN(s_logisimNet70),
.clock(s_logisimNet111),
.func(s_logisimBus58[5:0]),
.j(s_logisimNet55),
.jal(s_logisimNet50),
.jr(s_logisimNet57),
.link(s_logisimNet67),
.memToReg(s_logisimNet64),
.memWrite(s_logisimNet25),
.opCode(s_logisimBus22[5:0]),
.regDst(s_logisimNet45),
.regWrite(s_logisimNet60),
.rst(s_logisimNet77),
.shift(s_logisimNet26));
endmodule