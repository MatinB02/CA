/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
CU4
**
**
**
*****************************************************************************/
module
CU4(
memWrite,
opCode
);
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
[5:0]
opCode;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
memWrite;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
[5:0]
s_logisimBus1;
wire
[5:0]
s_logisimBus2;
wire
s_logisimNet0;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
all
input
connections
are
defined
**
*******************************************************************************/
assign
s_logisimBus1[5:0]
=
opCode;
/*******************************************************************************
**
Here
all
output
connections
are
defined
**
*******************************************************************************/
assign
memWrite
=
s_logisimNet0;
/*******************************************************************************
**
Here
all
in-lined
components
are
defined
**
*******************************************************************************/
assign
s_logisimBus2[5:0]
=
{2'b10,
4'hB};
/*******************************************************************************
**
Here
all
normal
components
are
defined
**
*******************************************************************************/
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_1
(.aEqualsB(s_logisimNet0),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus2[5:0]),
.dataB(s_logisimBus1[5:0]));
endmodule