/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
XORR
**
**
**
*****************************************************************************/
module
XORR(
a,
b,
res_high,
res_low
);
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
[31:0]
a;
input
[31:0]
b;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
[31:0]
res_high;
output
[31:0]
res_low;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
[31:0]
s_logisimBus0;
wire
[31:0]
s_logisimBus1;
wire
[31:0]
s_logisimBus2;
wire
[31:0]
s_logisimBus3;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
all
input
connections
are
defined
**
*******************************************************************************/
assign
s_logisimBus1[31:0]
=
a;
assign
s_logisimBus2[31:0]
=
b;
/*******************************************************************************
**
Here
all
output
connections
are
defined
**
*******************************************************************************/
assign
res_high
=
s_logisimBus0[31:0];
assign
res_low
=
s_logisimBus3[31:0];
/*******************************************************************************
**
Here
all
in-lined
components
are
defined
**
*******************************************************************************/
assign
s_logisimBus0[31:0]
=
32'h00000000;
/*******************************************************************************
**
Here
all
normal
components
are
defined
**
*******************************************************************************/
XOR_GATE_BUS_ONEHOT
#(.BubblesMask(2'b00),
.NrOfBits(32))
GATES_1
(.input1(s_logisimBus1[31:0]),
.input2(s_logisimBus2[31:0]),
.result(s_logisimBus3[31:0]));
endmodule