/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
InstructionDecode
**
**
**
*****************************************************************************/
module
InstructionDecode(
Instruction,
Itype,
func,
imm,
rd,
rs,
rt,
shmt
);
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
[31:0]
Instruction;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
Itype;
output
[5:0]
func;
output
[15:0]
imm;
output
[4:0]
rd;
output
[4:0]
rs;
output
[4:0]
rt;
output
[4:0]
shmt;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
[31:0]
s_logisimBus2;
wire
[5:0]
s_logisimBus9;
wire
s_logisimNet6;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
all
input
connections
are
defined
**
*******************************************************************************/
assign
s_logisimBus2[31:0]
=
Instruction;
/*******************************************************************************
**
Here
all
output
connections
are
defined
**
*******************************************************************************/
assign
Itype
=
s_logisimNet6;
assign
func
=
s_logisimBus2[5:0];
assign
imm
=
s_logisimBus2[15:0];
assign
rd
=
s_logisimBus2[15:11];
assign
rs
=
s_logisimBus2[20:16];
assign
rt
=
s_logisimBus2[25:21];
assign
shmt
=
s_logisimBus2[10:6];
/*******************************************************************************
**
Here
all
in-lined
components
are
defined
**
*******************************************************************************/
assign
s_logisimBus9[5:0]
=
{2'b00,
4'h0};
/*******************************************************************************
**
Here
all
normal
components
are
defined
**
*******************************************************************************/
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_1
(.aEqualsB(),
.aGreaterThanB(),
.aLessThanB(s_logisimNet6),
.dataA(s_logisimBus9[5:0]),
.dataB(s_logisimBus2[31:26]));
endmodule