/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
FAA
**
**
**
*****************************************************************************/
module
FAA(
a,
b,
c,
cout,
s
);
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
[63:0]
a;
input
[63:0]
b;
input
[63:0]
c;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
[63:0]
cout;
output
[63:0]
s;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
[63:0]
s_logisimBus0;
wire
[63:0]
s_logisimBus1;
wire
[63:0]
s_logisimBus2;
wire
[63:0]
s_logisimBus3;
wire
[63:0]
s_logisimBus4;
wire
[63:0]
s_logisimBus5;
wire
[63:0]
s_logisimBus6;
wire
[63:0]
s_logisimBus7;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
all
input
connections
are
defined
**
*******************************************************************************/
assign
s_logisimBus0[63:0]
=
a;
assign
s_logisimBus1[63:0]
=
c;
assign
s_logisimBus2[63:0]
=
b;
/*******************************************************************************
**
Here
all
output
connections
are
defined
**
*******************************************************************************/
assign
cout
=
s_logisimBus6[63:0];
assign
s
=
s_logisimBus5[63:0];
/*******************************************************************************
**
Here
all
normal
components
are
defined
**
*******************************************************************************/
AND_GATE_BUS
#(.BubblesMask(2'b00),
.NrOfBits(64))
GATES_1
(.input1(s_logisimBus2[63:0]),
.input2(s_logisimBus0[63:0]),
.result(s_logisimBus7[63:0]));
XOR_GATE_BUS_ONEHOT
#(.BubblesMask(2'b00),
.NrOfBits(64))
GATES_2
(.input1(s_logisimBus0[63:0]),
.input2(s_logisimBus2[63:0]),
.result(s_logisimBus4[63:0]));
AND_GATE_BUS
#(.BubblesMask(2'b00),
.NrOfBits(64))
GATES_3
(.input1(s_logisimBus4[63:0]),
.input2(s_logisimBus1[63:0]),
.result(s_logisimBus3[63:0]));
XOR_GATE_BUS_ONEHOT
#(.BubblesMask(2'b00),
.NrOfBits(64))
GATES_4
(.input1(s_logisimBus4[63:0]),
.input2(s_logisimBus1[63:0]),
.result(s_logisimBus5[63:0]));
OR_GATE_BUS
#(.BubblesMask(2'b00),
.NrOfBits(64))
GATES_5
(.input1(s_logisimBus7[63:0]),
.input2(s_logisimBus3[63:0]),
.result(s_logisimBus6[63:0]));
endmodule