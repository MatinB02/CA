/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
ROTRR
**
**
**
*****************************************************************************/
module
ROTRR(
a,
b,
res_high,
res_low
);
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
[31:0]
a;
input
[31:0]
b;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
[31:0]
res_high;
output
[31:0]
res_low;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
[31:0]
s_logisimBus0;
wire
[31:0]
s_logisimBus2;
wire
[63:0]
s_logisimBus5;
wire
[31:0]
s_logisimBus6;
wire
[63:0]
s_logisimBus8;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
all
input
connections
are
defined
**
*******************************************************************************/
assign
s_logisimBus2[31:0]
=
b;
assign
s_logisimBus5[63:32]
=
a;
/*******************************************************************************
**
Here
all
output
connections
are
defined
**
*******************************************************************************/
assign
res_high
=
s_logisimBus6[31:0];
assign
res_low
=
s_logisimBus0[31:0];
/*******************************************************************************
**
Here
all
in-lined
components
are
defined
**
*******************************************************************************/
assign
s_logisimBus5[31:0]
=
32'h00000000;
assign
s_logisimBus6[31:0]
=
32'h00000000;
/*******************************************************************************
**
Here
all
normal
components
are
defined
**
*******************************************************************************/
OR_GATE_BUS
#(.BubblesMask(2'b00),
.NrOfBits(32))
GATES_1
(.input1(s_logisimBus8[31:0]),
.input2(s_logisimBus8[63:32]),
.result(s_logisimBus0[31:0]));
/*******************************************************************************
**
Here
all
sub-circuits
are
defined
**
*******************************************************************************/
SRL64
SRL64_1
(.a(s_logisimBus5[63:0]),
.b(s_logisimBus2[31:0]),
.res_high(),
.res_low(s_logisimBus8[63:0]));
endmodule