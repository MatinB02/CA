/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
main
**
**
**
*****************************************************************************/
module
main(
a,
aluop,
b,
clk,
done,
output_inc,
output_inverted,
res_high,
res_low,
rst
);
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
[31:0]
a;
input
[3:0]
aluop;
input
[31:0]
b;
input
clk;
input
output_inc;
input
output_inverted;
input
rst;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
done;
output
[31:0]
res_high;
output
[31:0]
res_low;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
[31:0]
s_logisimBus0;
wire
[31:0]
s_logisimBus1;
wire
[31:0]
s_logisimBus10;
wire
[31:0]
s_logisimBus12;
wire
[63:0]
s_logisimBus13;
wire
[31:0]
s_logisimBus15;
wire
[31:0]
s_logisimBus16;
wire
[31:0]
s_logisimBus17;
wire
[31:0]
s_logisimBus19;
wire
[31:0]
s_logisimBus2;
wire
[31:0]
s_logisimBus21;
wire
[31:0]
s_logisimBus22;
wire
[31:0]
s_logisimBus23;
wire
[31:0]
s_logisimBus24;
wire
[31:0]
s_logisimBus25;
wire
[31:0]
s_logisimBus27;
wire
[31:0]
s_logisimBus28;
wire
[31:0]
s_logisimBus29;
wire
[31:0]
s_logisimBus3;
wire
[31:0]
s_logisimBus30;
wire
[63:0]
s_logisimBus31;
wire
[31:0]
s_logisimBus33;
wire
[31:0]
s_logisimBus34;
wire
[31:0]
s_logisimBus35;
wire
[31:0]
s_logisimBus36;
wire
[63:0]
s_logisimBus4;
wire
[63:0]
s_logisimBus40;
wire
[63:0]
s_logisimBus41;
wire
[63:0]
s_logisimBus42;
wire
[63:0]
s_logisimBus43;
wire
[3:0]
s_logisimBus44;
wire
[31:0]
s_logisimBus45;
wire
[31:0]
s_logisimBus5;
wire
[3:0]
s_logisimBus7;
wire
[31:0]
s_logisimBus8;
wire
[31:0]
s_logisimBus9;
wire
s_logisimNet14;
wire
s_logisimNet20;
wire
s_logisimNet26;
wire
s_logisimNet32;
wire
s_logisimNet37;
wire
s_logisimNet6;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
all
input
connections
are
defined
**
*******************************************************************************/
assign
s_logisimBus1[31:0]
=
a;
assign
s_logisimBus24[31:0]
=
b;
assign
s_logisimBus7[3:0]
=
aluop;
assign
s_logisimNet20
=
output_inc;
assign
s_logisimNet26
=
rst;
assign
s_logisimNet37
=
output_inverted;
assign
s_logisimNet6
=
clk;
/*******************************************************************************
**
Here
all
output
connections
are
defined
**
*******************************************************************************/
assign
done
=
s_logisimNet32;
assign
res_high
=
s_logisimBus13[63:32];
assign
res_low
=
s_logisimBus13[31:0];
/*******************************************************************************
**
Here
all
in-lined
components
are
defined
**
*******************************************************************************/
assign
s_logisimBus42[63:0]
=
64'h0000000000000001;
assign
s_logisimNet32
=
1'b1;
assign
s_logisimBus44[3:0]
=
4'h1;
assign
s_logisimBus43
=
~s_logisimBus31;
assign
s_logisimBus45
=
~s_logisimBus1;
/*******************************************************************************
**
Here
all
normal
components
are
defined
**
*******************************************************************************/
Multiplexer_bus_2
#(.nrOfBits(64))
PLEXERS_1
(.enable(1'b1),
.muxIn_0(s_logisimBus31[63:0]),
.muxIn_1(s_logisimBus43[63:0]),
.muxOut(s_logisimBus4[63:0]),
.sel(s_logisimNet37));
Multiplexer_bus_2
#(.nrOfBits(64))
PLEXERS_2
(.enable(1'b1),
.muxIn_0(s_logisimBus4[63:0]),
.muxIn_1(s_logisimBus40[63:0]),
.muxOut(s_logisimBus13[63:0]),
.sel(s_logisimNet20));
Multiplexer_bus_16
#(.nrOfBits(32))
PLEXERS_3
(.enable(1'b1),
.muxIn_0(s_logisimBus33[31:0]),
.muxIn_1(s_logisimBus33[31:0]),
.muxIn_10(s_logisimBus8[31:0]),
.muxIn_11(s_logisimBus19[31:0]),
.muxIn_12(s_logisimBus35[31:0]),
.muxIn_13(32'd0),
.muxIn_14(32'd0),
.muxIn_15(32'd0),
.muxIn_2(s_logisimBus12[31:0]),
.muxIn_3(s_logisimBus36[31:0]),
.muxIn_4(s_logisimBus2[31:0]),
.muxIn_5(s_logisimBus27[31:0]),
.muxIn_6(s_logisimBus34[31:0]),
.muxIn_7(s_logisimBus0[31:0]),
.muxIn_8(s_logisimBus30[31:0]),
.muxIn_9(s_logisimBus5[31:0]),
.muxOut(s_logisimBus41[63:32]),
.sel(s_logisimBus7[3:0]));
Multiplexer_bus_16
#(.nrOfBits(32))
PLEXERS_4
(.enable(1'b1),
.muxIn_0(s_logisimBus17[31:0]),
.muxIn_1(s_logisimBus17[31:0]),
.muxIn_10(s_logisimBus21[31:0]),
.muxIn_11(s_logisimBus22[31:0]),
.muxIn_12(s_logisimBus15[31:0]),
.muxIn_13(32'd0),
.muxIn_14(32'd0),
.muxIn_15(32'd0),
.muxIn_2(s_logisimBus25[31:0]),
.muxIn_3(s_logisimBus29[31:0]),
.muxIn_4(s_logisimBus3[31:0]),
.muxIn_5(s_logisimBus9[31:0]),
.muxIn_6(s_logisimBus28[31:0]),
.muxIn_7(s_logisimBus23[31:0]),
.muxIn_8(s_logisimBus10[31:0]),
.muxIn_9(s_logisimBus16[31:0]),
.muxOut(s_logisimBus41[31:0]),
.sel(s_logisimBus7[3:0]));
Adder
#(.extendedBits(65),
.nrOfBits(64))
ARITH_5
(.carryIn(1'b0),
.carryOut(),
.dataA(s_logisimBus4[63:0]),
.dataB(s_logisimBus42[63:0]),
.result(s_logisimBus40[63:0]));
Comparator
#(.nrOfBits(4),
.twosComplement(0))
ARITH_6
(.aEqualsB(s_logisimNet14),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus7[3:0]),
.dataB(s_logisimBus44[3:0]));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(64))
MEMORY_7
(.clock(s_logisimNet6),
.clockEnable(1'b1),
.d(s_logisimBus41[63:0]),
.q(s_logisimBus31[63:0]),
.reset(s_logisimNet26),
.tick(1'b1));
/*******************************************************************************
**
Here
all
sub-circuits
are
defined
**
*******************************************************************************/
CLOO
CLOO_1
(.a(s_logisimBus1[31:0]),
.res_high(s_logisimBus0[31:0]),
.res_low(s_logisimBus23[31:0]));
CLOO
CLOO_2
(.a(s_logisimBus45[31:0]),
.res_high(s_logisimBus30[31:0]),
.res_low(s_logisimBus10[31:0]));
MULL
MULL_1
(.Done(),
.a(s_logisimBus1[31:0]),
.b(s_logisimBus24[31:0]),
.clk(s_logisimNet6),
.res_high(s_logisimBus12[31:0]),
.res_low(s_logisimBus25[31:0]));
ADDD
ADDD_1
(.Output_bus_1(),
.S(s_logisimNet14),
.a(s_logisimBus1[31:0]),
.b(s_logisimBus24[31:0]),
.res_high(s_logisimBus33[31:0]),
.res_low(s_logisimBus17[31:0]));
DIVV
DIVV_1
(.clk(s_logisimNet6),
.dividend(s_logisimBus1[31:0]),
.divisor(s_logisimBus24[31:0]),
.done(),
.quotient(s_logisimBus29[31:0]),
.remainder(s_logisimBus36[31:0]));
ANDD
ANDD_1
(.a(s_logisimBus1[31:0]),
.b(s_logisimBus24[31:0]),
.res_high(s_logisimBus2[31:0]),
.res_low(s_logisimBus3[31:0]));
ORR
ORR_1
(.a(s_logisimBus1[31:0]),
.b(s_logisimBus24[31:0]),
.res_high(s_logisimBus27[31:0]),
.res_low(s_logisimBus9[31:0]));
XORR
XORR_1
(.a(s_logisimBus1[31:0]),
.b(s_logisimBus24[31:0]),
.res_high(s_logisimBus34[31:0]),
.res_low(s_logisimBus28[31:0]));
SLLL
SLLL_1
(.a(s_logisimBus1[31:0]),
.b(s_logisimBus24[31:0]),
.res_high(s_logisimBus5[31:0]),
.res_low(s_logisimBus16[31:0]));
SRLL
SRLL_1
(.a(s_logisimBus1[31:0]),
.b(s_logisimBus24[31:0]),
.res_high(s_logisimBus8[31:0]),
.res_low(s_logisimBus21[31:0]));
SRAA
SRAA_1
(.a(s_logisimBus1[31:0]),
.b(s_logisimBus24[31:0]),
.res_high(s_logisimBus19[31:0]),
.res_low(s_logisimBus22[31:0]));
ROTRR
ROTRR_1
(.a(s_logisimBus1[31:0]),
.b(s_logisimBus24[31:0]),
.res_high(s_logisimBus35[31:0]),
.res_low(s_logisimBus15[31:0]));
endmodule