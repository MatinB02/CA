/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
ControlUnit
**
**
**
*****************************************************************************/
module
ControlUnit(
ALUop,
ALUsrc,
FALUop,
FROMCOP,
FregWrite,
TOCOP,
branch,
divv,
first,
fsin,
func,
inst,
j,
main_clock,
memToReg,
memWrite,
mohi,
nop,
opCode,
pc,
regDst,
regWrite,
shmt
);
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
[5:0]
func;
input
inst;
input
main_clock;
input
[5:0]
opCode;
input
[8:0]
pc;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
[3:0]
ALUop;
output
ALUsrc;
output
[2:0]
FALUop;
output
FROMCOP;
output
FregWrite;
output
TOCOP;
output
branch;
output
divv;
output
first;
output
fsin;
output
j;
output
memToReg;
output
memWrite;
output
mohi;
output
nop;
output
regDst;
output
regWrite;
output
shmt;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
[5:0]
s_logisimBus10;
wire
[3:0]
s_logisimBus100;
wire
[3:0]
s_logisimBus101;
wire
[3:0]
s_logisimBus102;
wire
[3:0]
s_logisimBus103;
wire
[3:0]
s_logisimBus104;
wire
[5:0]
s_logisimBus105;
wire
[5:0]
s_logisimBus106;
wire
[5:0]
s_logisimBus107;
wire
[5:0]
s_logisimBus108;
wire
[5:0]
s_logisimBus109;
wire
[5:0]
s_logisimBus110;
wire
[5:0]
s_logisimBus111;
wire
[5:0]
s_logisimBus112;
wire
[5:0]
s_logisimBus113;
wire
[5:0]
s_logisimBus114;
wire
[5:0]
s_logisimBus115;
wire
[5:0]
s_logisimBus116;
wire
[5:0]
s_logisimBus117;
wire
[5:0]
s_logisimBus118;
wire
[5:0]
s_logisimBus119;
wire
[5:0]
s_logisimBus120;
wire
[5:0]
s_logisimBus121;
wire
[5:0]
s_logisimBus122;
wire
[5:0]
s_logisimBus123;
wire
[5:0]
s_logisimBus124;
wire
[5:0]
s_logisimBus125;
wire
[5:0]
s_logisimBus126;
wire
[5:0]
s_logisimBus127;
wire
[5:0]
s_logisimBus128;
wire
[5:0]
s_logisimBus129;
wire
[5:0]
s_logisimBus130;
wire
[5:0]
s_logisimBus131;
wire
[5:0]
s_logisimBus132;
wire
[8:0]
s_logisimBus14;
wire
[3:0]
s_logisimBus18;
wire
[5:0]
s_logisimBus19;
wire
[2:0]
s_logisimBus20;
wire
[3:0]
s_logisimBus21;
wire
[3:0]
s_logisimBus22;
wire
[3:0]
s_logisimBus24;
wire
[8:0]
s_logisimBus33;
wire
[3:0]
s_logisimBus34;
wire
[3:0]
s_logisimBus35;
wire
[3:0]
s_logisimBus37;
wire
[3:0]
s_logisimBus42;
wire
[3:0]
s_logisimBus43;
wire
[2:0]
s_logisimBus44;
wire
[2:0]
s_logisimBus45;
wire
[2:0]
s_logisimBus47;
wire
[3:0]
s_logisimBus48;
wire
[3:0]
s_logisimBus50;
wire
[2:0]
s_logisimBus53;
wire
[3:0]
s_logisimBus56;
wire
[3:0]
s_logisimBus58;
wire
[3:0]
s_logisimBus59;
wire
[3:0]
s_logisimBus6;
wire
[2:0]
s_logisimBus60;
wire
[3:0]
s_logisimBus66;
wire
[3:0]
s_logisimBus68;
wire
[3:0]
s_logisimBus7;
wire
[2:0]
s_logisimBus72;
wire
[2:0]
s_logisimBus75;
wire
[2:0]
s_logisimBus76;
wire
[2:0]
s_logisimBus77;
wire
[3:0]
s_logisimBus78;
wire
[3:0]
s_logisimBus79;
wire
[2:0]
s_logisimBus80;
wire
[3:0]
s_logisimBus81;
wire
[2:0]
s_logisimBus82;
wire
[3:0]
s_logisimBus83;
wire
[2:0]
s_logisimBus84;
wire
[3:0]
s_logisimBus86;
wire
[2:0]
s_logisimBus87;
wire
[3:0]
s_logisimBus88;
wire
[2:0]
s_logisimBus89;
wire
[3:0]
s_logisimBus9;
wire
[3:0]
s_logisimBus90;
wire
[3:0]
s_logisimBus92;
wire
[3:0]
s_logisimBus93;
wire
[3:0]
s_logisimBus94;
wire
[3:0]
s_logisimBus95;
wire
[3:0]
s_logisimBus96;
wire
[3:0]
s_logisimBus97;
wire
[3:0]
s_logisimBus98;
wire
[3:0]
s_logisimBus99;
wire
s_logisimNet0;
wire
s_logisimNet1;
wire
s_logisimNet11;
wire
s_logisimNet12;
wire
s_logisimNet13;
wire
s_logisimNet133;
wire
s_logisimNet15;
wire
s_logisimNet16;
wire
s_logisimNet17;
wire
s_logisimNet2;
wire
s_logisimNet23;
wire
s_logisimNet25;
wire
s_logisimNet26;
wire
s_logisimNet27;
wire
s_logisimNet28;
wire
s_logisimNet29;
wire
s_logisimNet3;
wire
s_logisimNet30;
wire
s_logisimNet31;
wire
s_logisimNet32;
wire
s_logisimNet36;
wire
s_logisimNet38;
wire
s_logisimNet39;
wire
s_logisimNet4;
wire
s_logisimNet40;
wire
s_logisimNet41;
wire
s_logisimNet46;
wire
s_logisimNet49;
wire
s_logisimNet5;
wire
s_logisimNet51;
wire
s_logisimNet52;
wire
s_logisimNet54;
wire
s_logisimNet55;
wire
s_logisimNet57;
wire
s_logisimNet61;
wire
s_logisimNet62;
wire
s_logisimNet63;
wire
s_logisimNet64;
wire
s_logisimNet65;
wire
s_logisimNet67;
wire
s_logisimNet69;
wire
s_logisimNet70;
wire
s_logisimNet71;
wire
s_logisimNet73;
wire
s_logisimNet74;
wire
s_logisimNet8;
wire
s_logisimNet85;
wire
s_logisimNet91;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
all
input
connections
are
defined
**
*******************************************************************************/
assign
s_logisimBus10[5:0]
=
func;
assign
s_logisimBus19[5:0]
=
opCode;
assign
s_logisimBus33[8:0]
=
pc;
assign
s_logisimNet13
=
inst;
assign
s_logisimNet133
=
main_clock;
/*******************************************************************************
**
Here
all
output
connections
are
defined
**
*******************************************************************************/
assign
ALUop
=
s_logisimBus66[3:0];
assign
ALUsrc
=
s_logisimNet74;
assign
FALUop
=
s_logisimBus47[2:0];
assign
FROMCOP
=
s_logisimNet63;
assign
FregWrite
=
s_logisimNet25;
assign
TOCOP
=
s_logisimNet57;
assign
branch
=
s_logisimNet69;
assign
divv
=
s_logisimNet26;
assign
first
=
s_logisimNet70;
assign
fsin
=
s_logisimNet15;
assign
j
=
s_logisimNet32;
assign
memToReg
=
s_logisimNet49;
assign
memWrite
=
s_logisimNet54;
assign
mohi
=
s_logisimNet29;
assign
nop
=
s_logisimNet31;
assign
regDst
=
s_logisimNet65;
assign
regWrite
=
s_logisimNet73;
assign
shmt
=
s_logisimNet12;
/*******************************************************************************
**
Here
all
in-lined
components
are
defined
**
*******************************************************************************/
assign
s_logisimBus107[5:0]
=
{2'b10,
4'h0};
assign
s_logisimBus105[5:0]
=
{2'b01,
4'h4};
assign
s_logisimBus106[5:0]
=
{2'b01,
4'h5};
assign
s_logisimBus108[5:0]
=
{2'b01,
4'h6};
assign
s_logisimBus109[5:0]
=
{2'b01,
4'h7};
assign
s_logisimBus110[5:0]
=
{2'b01,
4'h8};
assign
s_logisimBus111[5:0]
=
{2'b01,
4'h9};
assign
s_logisimBus112[5:0]
=
{2'b10,
4'h2};
assign
s_logisimBus113[5:0]
=
{2'b10,
4'h4};
assign
s_logisimBus114[5:0]
=
{2'b10,
4'h5};
assign
s_logisimBus115[5:0]
=
{2'b10,
4'h6};
assign
s_logisimBus116[5:0]
=
{2'b00,
4'h4};
assign
s_logisimBus117[5:0]
=
{2'b00,
4'h6};
assign
s_logisimBus118[5:0]
=
{2'b00,
4'h7};
assign
s_logisimBus119[5:0]
=
{2'b01,
4'hA};
assign
s_logisimBus120[5:0]
=
{2'b01,
4'h0};
assign
s_logisimBus121[5:0]
=
{2'b00,
4'h0};
assign
s_logisimBus122[5:0]
=
{2'b00,
4'h8};
assign
s_logisimBus123[5:0]
=
{2'b01,
4'h2};
assign
s_logisimBus124[5:0]
=
{2'b00,
4'h1};
assign
s_logisimBus125[5:0]
=
{2'b01,
4'h3};
assign
s_logisimBus75[2:0]
=
3'b111;
assign
s_logisimBus76[2:0]
=
3'b101;
assign
s_logisimBus77[2:0]
=
3'b100;
assign
s_logisimBus78[3:0]
=
4'hF;
assign
s_logisimBus79[3:0]
=
4'h0;
assign
s_logisimBus80[2:0]
=
3'b011;
assign
s_logisimBus81[3:0]
=
4'h1;
assign
s_logisimBus82[2:0]
=
3'b010;
assign
s_logisimBus83[3:0]
=
4'h4;
assign
s_logisimBus84[2:0]
=
3'b001;
assign
s_logisimNet85
=
1'b1;
assign
s_logisimBus86[3:0]
=
4'h5;
assign
s_logisimBus87[2:0]
=
3'b000;
assign
s_logisimBus88[3:0]
=
4'h6;
assign
s_logisimBus89[2:0]
=
3'b111;
assign
s_logisimBus90[3:0]
=
4'h9;
assign
s_logisimNet91
=
1'b0;
assign
s_logisimBus92[3:0]
=
4'hA;
assign
s_logisimBus93[3:0]
=
4'hB;
assign
s_logisimBus126[5:0]
=
{2'b00,
4'h0};
assign
s_logisimBus127[5:0]
=
{2'b00,
4'h8};
assign
s_logisimBus128[5:0]
=
{2'b10,
4'hB};
assign
s_logisimBus129[5:0]
=
{2'b10,
4'h3};
assign
s_logisimBus130[5:0]
=
{2'b00,
4'h5};
assign
s_logisimBus131[5:0]
=
{2'b00,
4'hA};
assign
s_logisimBus132[5:0]
=
{2'b00,
4'h2};
assign
s_logisimBus94[3:0]
=
4'h3;
assign
s_logisimBus95[3:0]
=
4'hF;
assign
s_logisimBus96[3:0]
=
4'h9;
assign
s_logisimBus97[3:0]
=
4'hF;
assign
s_logisimBus98[3:0]
=
4'hF;
assign
s_logisimBus99[3:0]
=
4'hC;
assign
s_logisimBus100[3:0]
=
4'h0;
assign
s_logisimBus101[3:0]
=
4'h0;
assign
s_logisimBus102[3:0]
=
4'h7;
assign
s_logisimBus103[3:0]
=
4'h2;
assign
s_logisimBus104[3:0]
=
4'hF;
assign
s_logisimNet71
=
~s_logisimNet13;
assign
s_logisimNet70
=
~s_logisimNet2;
/*******************************************************************************
**
Here
all
normal
components
are
defined
**
*******************************************************************************/
OR_GATE
#(.BubblesMask(2'b00))
GATES_1
(.input1(1'b0),
.input2(s_logisimNet39),
.result(s_logisimNet31));
OR_GATE_7_INPUTS
#(.BubblesMask({3'b000,
4'h0}))
GATES_2
(.input1(s_logisimNet61),
.input2(s_logisimNet38),
.input3(s_logisimNet55),
.input4(s_logisimNet62),
.input5(s_logisimNet52),
.input6(s_logisimNet40),
.input7(s_logisimNet57),
.result(s_logisimNet51));
AND_GATE
#(.BubblesMask(2'b00))
GATES_3
(.input1(s_logisimNet65),
.input2(s_logisimNet16),
.result(s_logisimNet29));
AND_GATE
#(.BubblesMask(2'b10))
GATES_4
(.input1(s_logisimNet13),
.input2(s_logisimNet23),
.result(s_logisimNet1));
AND_GATE
#(.BubblesMask(2'b00))
GATES_5
(.input1(s_logisimNet63),
.input2(s_logisimNet65),
.result(s_logisimNet5));
AND_GATE
#(.BubblesMask(2'b01))
GATES_6
(.input1(s_logisimNet51),
.input2(s_logisimNet65),
.result(s_logisimNet28));
AND_GATE
#(.BubblesMask(2'b00))
GATES_7
(.input1(s_logisimNet51),
.input2(s_logisimNet65),
.result(s_logisimNet25));
OR_GATE_5_INPUTS
#(.BubblesMask({1'b0,
4'h0}))
GATES_8
(.input1(s_logisimNet28),
.input2(s_logisimNet5),
.input3(s_logisimNet67),
.input4(s_logisimNet64),
.input5(s_logisimNet49),
.result(s_logisimNet73));
AND_GATE
#(.BubblesMask(2'b00))
GATES_9
(.input1(s_logisimNet61),
.input2(s_logisimNet65),
.result(s_logisimNet15));
OR_GATE_5_INPUTS
#(.BubblesMask({1'b0,
4'h0}))
GATES_10
(.input1(s_logisimNet67),
.input2(s_logisimNet54),
.input3(s_logisimNet49),
.input4(s_logisimNet69),
.input5(s_logisimNet64),
.result(s_logisimNet74));
Multiplexer_bus_2
#(.nrOfBits(3))
PLEXERS_11
(.enable(1'b1),
.muxIn_0(s_logisimBus75[2:0]),
.muxIn_1(s_logisimBus76[2:0]),
.muxOut(s_logisimBus44[2:0]),
.sel(s_logisimNet61));
Multiplexer_bus_2
#(.nrOfBits(3))
PLEXERS_12
(.enable(1'b1),
.muxIn_0(s_logisimBus44[2:0]),
.muxIn_1(s_logisimBus77[2:0]),
.muxOut(s_logisimBus60[2:0]),
.sel(s_logisimNet40));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_13
(.enable(1'b1),
.muxIn_0(s_logisimBus78[3:0]),
.muxIn_1(s_logisimBus79[3:0]),
.muxOut(s_logisimBus7[3:0]),
.sel(s_logisimNet3));
Multiplexer_bus_2
#(.nrOfBits(3))
PLEXERS_14
(.enable(1'b1),
.muxIn_0(s_logisimBus60[2:0]),
.muxIn_1(s_logisimBus80[2:0]),
.muxOut(s_logisimBus72[2:0]),
.sel(s_logisimNet52));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_15
(.enable(1'b1),
.muxIn_0(s_logisimBus7[3:0]),
.muxIn_1(s_logisimBus81[3:0]),
.muxOut(s_logisimBus48[3:0]),
.sel(s_logisimNet8));
Multiplexer_bus_2
#(.nrOfBits(3))
PLEXERS_16
(.enable(1'b1),
.muxIn_0(s_logisimBus72[2:0]),
.muxIn_1(s_logisimBus82[2:0]),
.muxOut(s_logisimBus20[2:0]),
.sel(s_logisimNet62));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_17
(.enable(1'b1),
.muxIn_0(s_logisimBus48[3:0]),
.muxIn_1(s_logisimBus83[3:0]),
.muxOut(s_logisimBus34[3:0]),
.sel(s_logisimNet41));
Multiplexer_bus_2
#(.nrOfBits(3))
PLEXERS_18
(.enable(1'b1),
.muxIn_0(s_logisimBus20[2:0]),
.muxIn_1(s_logisimBus84[2:0]),
.muxOut(s_logisimBus45[2:0]),
.sel(s_logisimNet55));
Multiplexer_2
PLEXERS_19
(.enable(1'b1),
.muxIn_0(s_logisimNet71),
.muxIn_1(s_logisimNet85),
.muxOut(s_logisimNet30),
.sel(s_logisimNet1));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_20
(.enable(1'b1),
.muxIn_0(s_logisimBus34[3:0]),
.muxIn_1(s_logisimBus86[3:0]),
.muxOut(s_logisimBus21[3:0]),
.sel(s_logisimNet4));
Multiplexer_bus_2
#(.nrOfBits(3))
PLEXERS_21
(.enable(1'b1),
.muxIn_0(s_logisimBus45[2:0]),
.muxIn_1(s_logisimBus87[2:0]),
.muxOut(s_logisimBus53[2:0]),
.sel(s_logisimNet38));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_22
(.enable(1'b1),
.muxIn_0(s_logisimBus21[3:0]),
.muxIn_1(s_logisimBus88[3:0]),
.muxOut(s_logisimBus6[3:0]),
.sel(s_logisimNet17));
Multiplexer_bus_2
#(.nrOfBits(3))
PLEXERS_23
(.enable(1'b1),
.muxIn_0(s_logisimBus89[2:0]),
.muxIn_1(s_logisimBus53[2:0]),
.muxOut(s_logisimBus47[2:0]),
.sel(s_logisimNet65));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_24
(.enable(1'b1),
.muxIn_0(s_logisimBus6[3:0]),
.muxIn_1(s_logisimBus90[3:0]),
.muxOut(s_logisimBus35[3:0]),
.sel(s_logisimNet0));
Multiplexer_2
PLEXERS_25
(.enable(1'b1),
.muxIn_0(s_logisimNet91),
.muxIn_1(s_logisimNet30),
.muxOut(s_logisimNet39),
.sel(s_logisimNet26));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_26
(.enable(1'b1),
.muxIn_0(s_logisimBus35[3:0]),
.muxIn_1(s_logisimBus92[3:0]),
.muxOut(s_logisimBus22[3:0]),
.sel(s_logisimNet46));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_27
(.enable(1'b1),
.muxIn_0(s_logisimBus22[3:0]),
.muxIn_1(s_logisimBus93[3:0]),
.muxOut(s_logisimBus9[3:0]),
.sel(s_logisimNet36));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_28
(.enable(1'b1),
.muxIn_0(s_logisimBus9[3:0]),
.muxIn_1(s_logisimBus94[3:0]),
.muxOut(s_logisimBus56[3:0]),
.sel(s_logisimNet26));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_29
(.enable(1'b1),
.muxIn_0(s_logisimBus56[3:0]),
.muxIn_1(s_logisimBus95[3:0]),
.muxOut(s_logisimBus50[3:0]),
.sel(s_logisimNet16));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_30
(.enable(1'b1),
.muxIn_0(s_logisimBus50[3:0]),
.muxIn_1(s_logisimBus96[3:0]),
.muxOut(s_logisimBus37[3:0]),
.sel(s_logisimNet12));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_31
(.enable(1'b1),
.muxIn_0(s_logisimBus37[3:0]),
.muxIn_1(s_logisimBus97[3:0]),
.muxOut(s_logisimBus24[3:0]),
.sel(s_logisimNet27));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_32
(.enable(1'b1),
.muxIn_0(s_logisimBus24[3:0]),
.muxIn_1(s_logisimBus98[3:0]),
.muxOut(s_logisimBus42[3:0]),
.sel(s_logisimNet11));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_33
(.enable(1'b1),
.muxIn_0(s_logisimBus42[3:0]),
.muxIn_1(s_logisimBus99[3:0]),
.muxOut(s_logisimBus58[3:0]),
.sel(s_logisimNet67));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_34
(.enable(1'b1),
.muxIn_0(s_logisimBus58[3:0]),
.muxIn_1(s_logisimBus100[3:0]),
.muxOut(s_logisimBus68[3:0]),
.sel(s_logisimNet54));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_35
(.enable(1'b1),
.muxIn_0(s_logisimBus68[3:0]),
.muxIn_1(s_logisimBus101[3:0]),
.muxOut(s_logisimBus18[3:0]),
.sel(s_logisimNet49));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_36
(.enable(1'b1),
.muxIn_0(s_logisimBus18[3:0]),
.muxIn_1(s_logisimBus102[3:0]),
.muxOut(s_logisimBus43[3:0]),
.sel(s_logisimNet69));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_37
(.enable(1'b1),
.muxIn_0(s_logisimBus43[3:0]),
.muxIn_1(s_logisimBus103[3:0]),
.muxOut(s_logisimBus59[3:0]),
.sel(s_logisimNet64));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_38
(.enable(1'b1),
.muxIn_0(s_logisimBus59[3:0]),
.muxIn_1(s_logisimBus104[3:0]),
.muxOut(s_logisimBus66[3:0]),
.sel(s_logisimNet32));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_39
(.aEqualsB(s_logisimNet55),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus105[5:0]),
.dataB(s_logisimBus10[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_40
(.aEqualsB(s_logisimNet62),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus106[5:0]),
.dataB(s_logisimBus10[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_41
(.aEqualsB(s_logisimNet3),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus107[5:0]),
.dataB(s_logisimBus10[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_42
(.aEqualsB(s_logisimNet52),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus108[5:0]),
.dataB(s_logisimBus10[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_43
(.aEqualsB(s_logisimNet40),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus109[5:0]),
.dataB(s_logisimBus10[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_44
(.aEqualsB(s_logisimNet57),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus110[5:0]),
.dataB(s_logisimBus10[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_45
(.aEqualsB(s_logisimNet63),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus111[5:0]),
.dataB(s_logisimBus10[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_46
(.aEqualsB(s_logisimNet8),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus112[5:0]),
.dataB(s_logisimBus10[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_47
(.aEqualsB(s_logisimNet41),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus113[5:0]),
.dataB(s_logisimBus10[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_48
(.aEqualsB(s_logisimNet4),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus114[5:0]),
.dataB(s_logisimBus10[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_49
(.aEqualsB(s_logisimNet17),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus115[5:0]),
.dataB(s_logisimBus10[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_50
(.aEqualsB(s_logisimNet0),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus116[5:0]),
.dataB(s_logisimBus10[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_51
(.aEqualsB(s_logisimNet46),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus117[5:0]),
.dataB(s_logisimBus10[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_52
(.aEqualsB(s_logisimNet36),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus118[5:0]),
.dataB(s_logisimBus10[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_53
(.aEqualsB(s_logisimNet26),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus119[5:0]),
.dataB(s_logisimBus10[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_54
(.aEqualsB(s_logisimNet16),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus120[5:0]),
.dataB(s_logisimBus10[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_55
(.aEqualsB(s_logisimNet12),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus121[5:0]),
.dataB(s_logisimBus10[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_56
(.aEqualsB(s_logisimNet27),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus122[5:0]),
.dataB(s_logisimBus10[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_57
(.aEqualsB(s_logisimNet11),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus123[5:0]),
.dataB(s_logisimBus10[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_58
(.aEqualsB(s_logisimNet61),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus124[5:0]),
.dataB(s_logisimBus10[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_59
(.aEqualsB(s_logisimNet38),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus125[5:0]),
.dataB(s_logisimBus10[5:0]));
Comparator
#(.nrOfBits(9),
.twosComplement(0))
ARITH_60
(.aEqualsB(s_logisimNet2),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus33[8:0]),
.dataB(s_logisimBus14[8:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_61
(.aEqualsB(s_logisimNet65),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus126[5:0]),
.dataB(s_logisimBus19[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_62
(.aEqualsB(s_logisimNet67),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus127[5:0]),
.dataB(s_logisimBus19[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_63
(.aEqualsB(s_logisimNet54),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus128[5:0]),
.dataB(s_logisimBus19[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_64
(.aEqualsB(s_logisimNet49),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus129[5:0]),
.dataB(s_logisimBus19[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_65
(.aEqualsB(s_logisimNet69),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus130[5:0]),
.dataB(s_logisimBus19[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_66
(.aEqualsB(s_logisimNet64),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus131[5:0]),
.dataB(s_logisimBus19[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_67
(.aEqualsB(s_logisimNet32),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus132[5:0]),
.dataB(s_logisimBus19[5:0]));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(1))
MEMORY_68
(.clock(s_logisimNet133),
.clockEnable(1'b1),
.d(s_logisimNet13),
.q(s_logisimNet23),
.reset(1'b0),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(9))
MEMORY_69
(.clock(s_logisimNet133),
.clockEnable(1'b1),
.d(s_logisimBus33[8:0]),
.q(s_logisimBus14[8:0]),
.reset(1'b0),
.tick(1'b1));
endmodule