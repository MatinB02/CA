/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
fsinn
**
**
**
*****************************************************************************/
module
fsinn(
a,
b,
clk,
done,
fsin,
res
);
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
[31:0]
a;
input
[31:0]
b;
input
clk;
input
fsin;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
done;
output
[31:0]
res;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
[31:0]
s_logisimBus0;
wire
[4:0]
s_logisimBus10;
wire
[31:0]
s_logisimBus12;
wire
[4:0]
s_logisimBus13;
wire
[4:0]
s_logisimBus14;
wire
[31:0]
s_logisimBus15;
wire
[31:0]
s_logisimBus16;
wire
[31:0]
s_logisimBus17;
wire
[31:0]
s_logisimBus18;
wire
[31:0]
s_logisimBus19;
wire
[31:0]
s_logisimBus2;
wire
[31:0]
s_logisimBus20;
wire
[31:0]
s_logisimBus21;
wire
[31:0]
s_logisimBus22;
wire
[31:0]
s_logisimBus23;
wire
[31:0]
s_logisimBus24;
wire
[31:0]
s_logisimBus25;
wire
[4:0]
s_logisimBus26;
wire
[31:0]
s_logisimBus27;
wire
[31:0]
s_logisimBus28;
wire
[31:0]
s_logisimBus29;
wire
[31:0]
s_logisimBus3;
wire
[31:0]
s_logisimBus30;
wire
[31:0]
s_logisimBus31;
wire
[31:0]
s_logisimBus32;
wire
[31:0]
s_logisimBus33;
wire
[31:0]
s_logisimBus34;
wire
[31:0]
s_logisimBus35;
wire
[31:0]
s_logisimBus36;
wire
[31:0]
s_logisimBus37;
wire
[31:0]
s_logisimBus38;
wire
[4:0]
s_logisimBus39;
wire
[4:0]
s_logisimBus4;
wire
[4:0]
s_logisimBus40;
wire
[31:0]
s_logisimBus41;
wire
[31:0]
s_logisimBus5;
wire
[4:0]
s_logisimBus6;
wire
[31:0]
s_logisimBus7;
wire
[31:0]
s_logisimBus8;
wire
s_logisimNet1;
wire
s_logisimNet11;
wire
s_logisimNet43;
wire
s_logisimNet9;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
all
input
connections
are
defined
**
*******************************************************************************/
assign
s_logisimBus25[31:0]
=
a;
assign
s_logisimBus3[31:0]
=
b;
assign
s_logisimNet11
=
fsin;
assign
s_logisimNet43
=
clk;
/*******************************************************************************
**
Here
all
output
connections
are
defined
**
*******************************************************************************/
assign
done
=
s_logisimNet9;
assign
res
=
s_logisimBus8[31:0];
/*******************************************************************************
**
Here
all
in-lined
components
are
defined
**
*******************************************************************************/
assign
s_logisimBus16[31:0]
=
32'h3F800000;
assign
s_logisimBus17[31:0]
=
32'h3C088889;
assign
s_logisimBus18[31:0]
=
32'h3638EF1D;
assign
s_logisimBus15[31:0]
=
32'h2F309231;
assign
s_logisimBus19[31:0]
=
32'h274A963C;
assign
s_logisimBus20[31:0]
=
32'h1EB8DC78;
assign
s_logisimBus21[31:0]
=
32'h159F9E67;
assign
s_logisimBus22[31:0]
=
32'h0C12CFCC;
assign
s_logisimBus23[31:0]
=
32'h021CC093;
assign
s_logisimBus24[31:0]
=
32'h00000034;
assign
s_logisimBus30[31:0]
=
32'hBE2AAAAB;
assign
s_logisimBus31[31:0]
=
32'hB9500D01;
assign
s_logisimBus29[31:0]
=
32'hB2D7322B;
assign
s_logisimBus28[31:0]
=
32'hAB573F9F;
assign
s_logisimBus27[31:0]
=
32'hA317A4DA;
assign
s_logisimBus32[31:0]
=
32'h9A3B0DA1;
assign
s_logisimBus33[31:0]
=
32'h90E8D58E;
assign
s_logisimBus34[31:0]
=
32'h8721A697;
assign
s_logisimBus35[31:0]
=
32'h80010DC6;
assign
s_logisimBus0[31:0]
=
32'h80000000;
assign
s_logisimBus5[31:0]
=
32'h0000001F;
assign
s_logisimBus6[4:0]
=
{1'b1,
4'hF};
assign
s_logisimBus39[4:0]
=
{1'b0,
4'h0};
assign
s_logisimBus40[4:0]
=
{1'b0,
4'h1};
/*******************************************************************************
**
Here
all
normal
components
are
defined
**
*******************************************************************************/
Multiplexer_bus_2
#(.nrOfBits(32))
PLEXERS_1
(.enable(1'b1),
.muxIn_0(s_logisimBus37[31:0]),
.muxIn_1(s_logisimBus25[31:0]),
.muxOut(s_logisimBus2[31:0]),
.sel(s_logisimNet11));
Multiplexer_bus_32
#(.nrOfBits(32))
PLEXERS_2
(.enable(1'b1),
.muxIn_0(s_logisimBus16[31:0]),
.muxIn_1(s_logisimBus30[31:0]),
.muxIn_10(s_logisimBus20[31:0]),
.muxIn_11(s_logisimBus32[31:0]),
.muxIn_12(s_logisimBus21[31:0]),
.muxIn_13(s_logisimBus33[31:0]),
.muxIn_14(s_logisimBus22[31:0]),
.muxIn_15(s_logisimBus34[31:0]),
.muxIn_16(s_logisimBus23[31:0]),
.muxIn_17(s_logisimBus35[31:0]),
.muxIn_18(s_logisimBus24[31:0]),
.muxIn_19(s_logisimBus0[31:0]),
.muxIn_2(s_logisimBus17[31:0]),
.muxIn_20(s_logisimBus0[31:0]),
.muxIn_21(s_logisimBus0[31:0]),
.muxIn_22(s_logisimBus0[31:0]),
.muxIn_23(s_logisimBus0[31:0]),
.muxIn_24(s_logisimBus0[31:0]),
.muxIn_25(s_logisimBus0[31:0]),
.muxIn_26(s_logisimBus0[31:0]),
.muxIn_27(s_logisimBus0[31:0]),
.muxIn_28(s_logisimBus0[31:0]),
.muxIn_29(s_logisimBus0[31:0]),
.muxIn_3(s_logisimBus31[31:0]),
.muxIn_30(s_logisimBus0[31:0]),
.muxIn_31(s_logisimBus0[31:0]),
.muxIn_4(s_logisimBus18[31:0]),
.muxIn_5(s_logisimBus29[31:0]),
.muxIn_6(s_logisimBus15[31:0]),
.muxIn_7(s_logisimBus28[31:0]),
.muxIn_8(s_logisimBus19[31:0]),
.muxIn_9(s_logisimBus27[31:0]),
.muxOut(s_logisimBus36[31:0]),
.sel(s_logisimBus4[4:0]));
Multiplexer_bus_2
#(.nrOfBits(5))
PLEXERS_3
(.enable(1'b1),
.muxIn_0(s_logisimBus3[4:0]),
.muxIn_1(s_logisimBus6[4:0]),
.muxOut(s_logisimBus13[4:0]),
.sel(s_logisimNet1));
Multiplexer_bus_2
#(.nrOfBits(5))
PLEXERS_4
(.enable(1'b1),
.muxIn_0(s_logisimBus10[4:0]),
.muxIn_1(s_logisimBus13[4:0]),
.muxOut(s_logisimBus14[4:0]),
.sel(s_logisimNet11));
Subtractor
#(.extendedBits(6),
.nrOfBits(5))
ARITH_5
(.borrowIn(1'b0),
.borrowOut(),
.dataA(s_logisimBus13[4:0]),
.dataB(s_logisimBus26[4:0]),
.result(s_logisimBus4[4:0]));
Comparator
#(.nrOfBits(32),
.twosComplement(0))
ARITH_6
(.aEqualsB(),
.aGreaterThanB(),
.aLessThanB(s_logisimNet1),
.dataA(s_logisimBus5[31:0]),
.dataB(s_logisimBus3[31:0]));
Comparator
#(.nrOfBits(5),
.twosComplement(0))
ARITH_7
(.aEqualsB(s_logisimNet9),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus26[4:0]),
.dataB(s_logisimBus39[4:0]));
Subtractor
#(.extendedBits(6),
.nrOfBits(5))
ARITH_8
(.borrowIn(1'b0),
.borrowOut(),
.dataA(s_logisimBus26[4:0]),
.dataB(s_logisimBus40[4:0]),
.result(s_logisimBus10[4:0]));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(32))
sum
(.clock(s_logisimNet43),
.clockEnable(1'b1),
.d(s_logisimBus12[31:0]),
.q(s_logisimBus8[31:0]),
.reset(s_logisimNet11),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(32))
x_powered
(.clock(s_logisimNet43),
.clockEnable(1'b1),
.d(s_logisimBus2[31:0]),
.q(s_logisimBus41[31:0]),
.reset(1'b0),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(5))
steps
(.clock(s_logisimNet43),
.clockEnable(1'b1),
.d(s_logisimBus14[4:0]),
.q(s_logisimBus26[4:0]),
.reset(1'b0),
.tick(1'b1));
/*******************************************************************************
**
Here
all
sub-circuits
are
defined
**
*******************************************************************************/
fadd
addh
(.INFINITY_PIN(),
.NAN_PIN(),
.a(s_logisimBus8[31:0]),
.b(s_logisimBus38[31:0]),
.res(s_logisimBus12[31:0]));
fmult
fmult_2
(.a(s_logisimBus41[31:0]),
.b(s_logisimBus7[31:0]),
.res(s_logisimBus37[31:0]));
fmult
multh
(.a(s_logisimBus41[31:0]),
.b(s_logisimBus36[31:0]),
.res(s_logisimBus38[31:0]));
fmult
fmult_1
(.a(s_logisimBus25[31:0]),
.b(s_logisimBus25[31:0]),
.res(s_logisimBus7[31:0]));
endmodule