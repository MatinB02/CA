/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
ControlUnit
**
**
**
*****************************************************************************/
module
ControlUnit(
ALUop,
ALUsrc,
Rtype,
beq,
branch,
divv,
func,
inst,
j,
jal,
jr,
main_clock,
memRead,
memToReg,
memWrite,
mohi,
mull,
nop,
opCode,
regDst,
regWrite,
shmt
);
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
[5:0]
func;
input
inst;
input
main_clock;
input
[5:0]
opCode;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
[3:0]
ALUop;
output
ALUsrc;
output
Rtype;
output
beq;
output
branch;
output
divv;
output
j;
output
jal;
output
jr;
output
memRead;
output
memToReg;
output
memWrite;
output
mohi;
output
mull;
output
nop;
output
regDst;
output
regWrite;
output
shmt;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
[5:0]
s_logisimBus10;
wire
[5:0]
s_logisimBus100;
wire
[5:0]
s_logisimBus101;
wire
[5:0]
s_logisimBus102;
wire
[5:0]
s_logisimBus103;
wire
[5:0]
s_logisimBus104;
wire
[5:0]
s_logisimBus105;
wire
[5:0]
s_logisimBus14;
wire
[3:0]
s_logisimBus15;
wire
[3:0]
s_logisimBus17;
wire
[3:0]
s_logisimBus18;
wire
[3:0]
s_logisimBus19;
wire
[3:0]
s_logisimBus2;
wire
[3:0]
s_logisimBus21;
wire
[3:0]
s_logisimBus22;
wire
[3:0]
s_logisimBus24;
wire
[3:0]
s_logisimBus26;
wire
[3:0]
s_logisimBus3;
wire
[3:0]
s_logisimBus32;
wire
[3:0]
s_logisimBus33;
wire
[3:0]
s_logisimBus35;
wire
[3:0]
s_logisimBus37;
wire
[3:0]
s_logisimBus39;
wire
[3:0]
s_logisimBus40;
wire
[3:0]
s_logisimBus45;
wire
[3:0]
s_logisimBus48;
wire
[3:0]
s_logisimBus5;
wire
[3:0]
s_logisimBus58;
wire
[3:0]
s_logisimBus59;
wire
[3:0]
s_logisimBus61;
wire
[3:0]
s_logisimBus62;
wire
[3:0]
s_logisimBus64;
wire
[3:0]
s_logisimBus65;
wire
[3:0]
s_logisimBus66;
wire
[3:0]
s_logisimBus67;
wire
[3:0]
s_logisimBus68;
wire
[3:0]
s_logisimBus69;
wire
[3:0]
s_logisimBus70;
wire
[3:0]
s_logisimBus71;
wire
[3:0]
s_logisimBus72;
wire
[3:0]
s_logisimBus73;
wire
[3:0]
s_logisimBus74;
wire
[3:0]
s_logisimBus75;
wire
[3:0]
s_logisimBus76;
wire
[3:0]
s_logisimBus77;
wire
[3:0]
s_logisimBus78;
wire
[3:0]
s_logisimBus79;
wire
[3:0]
s_logisimBus8;
wire
[3:0]
s_logisimBus80;
wire
[5:0]
s_logisimBus81;
wire
[5:0]
s_logisimBus82;
wire
[5:0]
s_logisimBus83;
wire
[5:0]
s_logisimBus84;
wire
[5:0]
s_logisimBus86;
wire
[5:0]
s_logisimBus87;
wire
[5:0]
s_logisimBus88;
wire
[5:0]
s_logisimBus89;
wire
[5:0]
s_logisimBus90;
wire
[5:0]
s_logisimBus91;
wire
[5:0]
s_logisimBus92;
wire
[5:0]
s_logisimBus93;
wire
[5:0]
s_logisimBus94;
wire
[5:0]
s_logisimBus95;
wire
[5:0]
s_logisimBus96;
wire
[5:0]
s_logisimBus97;
wire
[5:0]
s_logisimBus98;
wire
[5:0]
s_logisimBus99;
wire
s_logisimNet0;
wire
s_logisimNet1;
wire
s_logisimNet11;
wire
s_logisimNet12;
wire
s_logisimNet13;
wire
s_logisimNet16;
wire
s_logisimNet20;
wire
s_logisimNet23;
wire
s_logisimNet25;
wire
s_logisimNet27;
wire
s_logisimNet28;
wire
s_logisimNet29;
wire
s_logisimNet30;
wire
s_logisimNet31;
wire
s_logisimNet34;
wire
s_logisimNet36;
wire
s_logisimNet38;
wire
s_logisimNet4;
wire
s_logisimNet41;
wire
s_logisimNet42;
wire
s_logisimNet43;
wire
s_logisimNet44;
wire
s_logisimNet46;
wire
s_logisimNet47;
wire
s_logisimNet49;
wire
s_logisimNet50;
wire
s_logisimNet51;
wire
s_logisimNet52;
wire
s_logisimNet53;
wire
s_logisimNet54;
wire
s_logisimNet55;
wire
s_logisimNet56;
wire
s_logisimNet57;
wire
s_logisimNet6;
wire
s_logisimNet60;
wire
s_logisimNet63;
wire
s_logisimNet7;
wire
s_logisimNet85;
wire
s_logisimNet9;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
all
input
connections
are
defined
**
*******************************************************************************/
assign
s_logisimBus10[5:0]
=
func;
assign
s_logisimBus14[5:0]
=
opCode;
assign
s_logisimNet0
=
inst;
assign
s_logisimNet34
=
main_clock;
/*******************************************************************************
**
Here
all
output
connections
are
defined
**
*******************************************************************************/
assign
ALUop
=
s_logisimBus33[3:0];
assign
ALUsrc
=
s_logisimNet53;
assign
Rtype
=
s_logisimNet31;
assign
beq
=
s_logisimNet16;
assign
branch
=
s_logisimNet25;
assign
divv
=
s_logisimNet43;
assign
j
=
s_logisimNet36;
assign
jal
=
s_logisimNet20;
assign
jr
=
s_logisimNet44;
assign
memRead
=
s_logisimNet28;
assign
memToReg
=
s_logisimNet28;
assign
memWrite
=
s_logisimNet52;
assign
mohi
=
s_logisimNet41;
assign
mull
=
s_logisimNet57;
assign
nop
=
s_logisimNet29;
assign
regDst
=
s_logisimNet56;
assign
regWrite
=
s_logisimNet51;
assign
shmt
=
s_logisimNet38;
/*******************************************************************************
**
Here
all
in-lined
components
are
defined
**
*******************************************************************************/
assign
s_logisimBus81[5:0]
=
{2'b10,
4'h4};
assign
s_logisimBus84[5:0]
=
{2'b10,
4'h0};
assign
s_logisimBus82[5:0]
=
{2'b10,
4'h5};
assign
s_logisimBus83[5:0]
=
{2'b10,
4'h6};
assign
s_logisimBus86[5:0]
=
{2'b00,
4'h4};
assign
s_logisimBus87[5:0]
=
{2'b00,
4'h6};
assign
s_logisimBus88[5:0]
=
{2'b00,
4'h7};
assign
s_logisimBus89[5:0]
=
{2'b01,
4'hA};
assign
s_logisimBus90[5:0]
=
{2'b01,
4'h0};
assign
s_logisimBus91[5:0]
=
{2'b00,
4'h0};
assign
s_logisimBus92[5:0]
=
{2'b00,
4'h8};
assign
s_logisimBus93[5:0]
=
{2'b01,
4'h2};
assign
s_logisimBus95[5:0]
=
{2'b10,
4'h2};
assign
s_logisimBus94[5:0]
=
{2'b00,
4'h2};
assign
s_logisimBus58[3:0]
=
4'h0;
assign
s_logisimNet60
=
1'b1;
assign
s_logisimBus59[3:0]
=
4'h1;
assign
s_logisimBus61[3:0]
=
4'h4;
assign
s_logisimBus62[3:0]
=
4'h5;
assign
s_logisimNet63
=
1'b0;
assign
s_logisimBus64[3:0]
=
4'h6;
assign
s_logisimBus65[3:0]
=
4'h9;
assign
s_logisimBus96[5:0]
=
{2'b00,
4'h0};
assign
s_logisimBus97[5:0]
=
{2'b00,
4'h8};
assign
s_logisimBus98[5:0]
=
{2'b10,
4'hB};
assign
s_logisimBus99[5:0]
=
{2'b10,
4'h3};
assign
s_logisimBus100[5:0]
=
{2'b00,
4'h5};
assign
s_logisimBus101[5:0]
=
{2'b00,
4'hA};
assign
s_logisimBus102[5:0]
=
{2'b00,
4'h2};
assign
s_logisimBus103[5:0]
=
{2'b00,
4'h3};
assign
s_logisimBus104[5:0]
=
{2'b00,
4'h4};
assign
s_logisimBus105[5:0]
=
{2'b01,
4'hC};
assign
s_logisimBus66[3:0]
=
4'hA;
assign
s_logisimBus67[3:0]
=
4'hB;
assign
s_logisimBus68[3:0]
=
4'h3;
assign
s_logisimBus69[3:0]
=
4'hF;
assign
s_logisimBus70[3:0]
=
4'h9;
assign
s_logisimBus71[3:0]
=
4'hF;
assign
s_logisimBus72[3:0]
=
4'hF;
assign
s_logisimBus73[3:0]
=
4'hC;
assign
s_logisimBus74[3:0]
=
4'h0;
assign
s_logisimBus75[3:0]
=
4'h0;
assign
s_logisimBus76[3:0]
=
4'h7;
assign
s_logisimBus77[3:0]
=
4'h2;
assign
s_logisimBus78[3:0]
=
4'hF;
assign
s_logisimBus79[3:0]
=
4'h1;
assign
s_logisimBus80[3:0]
=
4'h8;
assign
s_logisimNet49
=
~s_logisimNet0;
/*******************************************************************************
**
Here
all
normal
components
are
defined
**
*******************************************************************************/
OR_GATE_5_INPUTS
#(.BubblesMask({1'b0,
4'h0}))
GATES_1
(.input1(s_logisimNet46),
.input2(s_logisimNet52),
.input3(s_logisimNet28),
.input4(s_logisimNet25),
.input5(s_logisimNet47),
.result(s_logisimNet53));
AND_GATE
#(.BubblesMask(2'b00))
GATES_2
(.input1(s_logisimNet44),
.input2(s_logisimNet31),
.result(s_logisimNet13));
OR_GATE_5_INPUTS
#(.BubblesMask({1'b0,
4'h0}))
GATES_3
(.input1(s_logisimNet13),
.input2(s_logisimNet46),
.input3(s_logisimNet57),
.input4(s_logisimNet47),
.input5(s_logisimNet28),
.result(s_logisimNet51));
AND_GATE
#(.BubblesMask(2'b00))
GATES_4
(.input1(s_logisimNet31),
.input2(s_logisimNet54),
.result(s_logisimNet41));
AND_GATE
#(.BubblesMask(2'b10))
GATES_5
(.input1(s_logisimNet0),
.input2(s_logisimNet7),
.result(s_logisimNet50));
AND_GATE
#(.BubblesMask(2'b00))
GATES_6
(.input1(s_logisimNet42),
.input2(s_logisimNet55),
.result(s_logisimNet57));
OR_GATE
#(.BubblesMask(2'b00))
GATES_7
(.input1(s_logisimNet57),
.input2(s_logisimNet31),
.result(s_logisimNet56));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_8
(.enable(1'b1),
.muxIn_0(s_logisimBus58[3:0]),
.muxIn_1(s_logisimBus59[3:0]),
.muxOut(s_logisimBus32[3:0]),
.sel(s_logisimNet6));
Multiplexer_2
PLEXERS_9
(.enable(1'b1),
.muxIn_0(s_logisimNet49),
.muxIn_1(s_logisimNet60),
.muxOut(s_logisimNet11),
.sel(s_logisimNet50));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_10
(.enable(1'b1),
.muxIn_0(s_logisimBus32[3:0]),
.muxIn_1(s_logisimBus61[3:0]),
.muxOut(s_logisimBus21[3:0]),
.sel(s_logisimNet27));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_11
(.enable(1'b1),
.muxIn_0(s_logisimBus21[3:0]),
.muxIn_1(s_logisimBus62[3:0]),
.muxOut(s_logisimBus15[3:0]),
.sel(s_logisimNet4));
Multiplexer_2
PLEXERS_12
(.enable(1'b1),
.muxIn_0(s_logisimNet63),
.muxIn_1(s_logisimNet11),
.muxOut(s_logisimNet29),
.sel(s_logisimNet43));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_13
(.enable(1'b1),
.muxIn_0(s_logisimBus15[3:0]),
.muxIn_1(s_logisimBus64[3:0]),
.muxOut(s_logisimBus5[3:0]),
.sel(s_logisimNet12));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_14
(.enable(1'b1),
.muxIn_0(s_logisimBus5[3:0]),
.muxIn_1(s_logisimBus65[3:0]),
.muxOut(s_logisimBus22[3:0]),
.sel(s_logisimNet1));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_15
(.enable(1'b1),
.muxIn_0(s_logisimBus22[3:0]),
.muxIn_1(s_logisimBus66[3:0]),
.muxOut(s_logisimBus17[3:0]),
.sel(s_logisimNet30));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_16
(.enable(1'b1),
.muxIn_0(s_logisimBus17[3:0]),
.muxIn_1(s_logisimBus67[3:0]),
.muxOut(s_logisimBus8[3:0]),
.sel(s_logisimNet23));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_17
(.enable(1'b1),
.muxIn_0(s_logisimBus8[3:0]),
.muxIn_1(s_logisimBus68[3:0]),
.muxOut(s_logisimBus40[3:0]),
.sel(s_logisimNet43));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_18
(.enable(1'b1),
.muxIn_0(s_logisimBus40[3:0]),
.muxIn_1(s_logisimBus69[3:0]),
.muxOut(s_logisimBus35[3:0]),
.sel(s_logisimNet54));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_19
(.enable(1'b1),
.muxIn_0(s_logisimBus35[3:0]),
.muxIn_1(s_logisimBus70[3:0]),
.muxOut(s_logisimBus26[3:0]),
.sel(s_logisimNet38));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_20
(.enable(1'b1),
.muxIn_0(s_logisimBus26[3:0]),
.muxIn_1(s_logisimBus71[3:0]),
.muxOut(s_logisimBus37[3:0]),
.sel(s_logisimNet44));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_21
(.enable(1'b1),
.muxIn_0(s_logisimBus37[3:0]),
.muxIn_1(s_logisimBus72[3:0]),
.muxOut(s_logisimBus45[3:0]),
.sel(s_logisimNet9));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_22
(.enable(1'b1),
.muxIn_0(s_logisimBus45[3:0]),
.muxIn_1(s_logisimBus73[3:0]),
.muxOut(s_logisimBus2[3:0]),
.sel(s_logisimNet46));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_23
(.enable(1'b1),
.muxIn_0(s_logisimBus2[3:0]),
.muxIn_1(s_logisimBus74[3:0]),
.muxOut(s_logisimBus19[3:0]),
.sel(s_logisimNet52));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_24
(.enable(1'b1),
.muxIn_0(s_logisimBus19[3:0]),
.muxIn_1(s_logisimBus75[3:0]),
.muxOut(s_logisimBus39[3:0]),
.sel(s_logisimNet28));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_25
(.enable(1'b1),
.muxIn_0(s_logisimBus39[3:0]),
.muxIn_1(s_logisimBus76[3:0]),
.muxOut(s_logisimBus48[3:0]),
.sel(s_logisimNet25));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_26
(.enable(1'b1),
.muxIn_0(s_logisimBus48[3:0]),
.muxIn_1(s_logisimBus77[3:0]),
.muxOut(s_logisimBus3[3:0]),
.sel(s_logisimNet47));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_27
(.enable(1'b1),
.muxIn_0(s_logisimBus3[3:0]),
.muxIn_1(s_logisimBus78[3:0]),
.muxOut(s_logisimBus18[3:0]),
.sel(s_logisimNet36));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_28
(.enable(1'b1),
.muxIn_0(s_logisimBus18[3:0]),
.muxIn_1(s_logisimBus79[3:0]),
.muxOut(s_logisimBus24[3:0]),
.sel(s_logisimNet16));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_29
(.enable(1'b1),
.muxIn_0(s_logisimBus24[3:0]),
.muxIn_1(s_logisimBus80[3:0]),
.muxOut(s_logisimBus33[3:0]),
.sel(s_logisimNet57));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_30
(.aEqualsB(s_logisimNet27),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus81[5:0]),
.dataB(s_logisimBus10[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_31
(.aEqualsB(s_logisimNet4),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus82[5:0]),
.dataB(s_logisimBus10[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_32
(.aEqualsB(s_logisimNet12),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus83[5:0]),
.dataB(s_logisimBus10[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_33
(.aEqualsB(s_logisimNet85),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus84[5:0]),
.dataB(s_logisimBus10[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_34
(.aEqualsB(s_logisimNet1),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus86[5:0]),
.dataB(s_logisimBus10[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_35
(.aEqualsB(s_logisimNet30),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus87[5:0]),
.dataB(s_logisimBus10[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_36
(.aEqualsB(s_logisimNet23),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus88[5:0]),
.dataB(s_logisimBus10[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_37
(.aEqualsB(s_logisimNet43),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus89[5:0]),
.dataB(s_logisimBus10[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_38
(.aEqualsB(s_logisimNet54),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus90[5:0]),
.dataB(s_logisimBus10[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_39
(.aEqualsB(s_logisimNet38),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus91[5:0]),
.dataB(s_logisimBus10[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_40
(.aEqualsB(s_logisimNet44),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus92[5:0]),
.dataB(s_logisimBus10[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_41
(.aEqualsB(s_logisimNet9),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus93[5:0]),
.dataB(s_logisimBus10[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_42
(.aEqualsB(s_logisimNet55),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus94[5:0]),
.dataB(s_logisimBus10[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_43
(.aEqualsB(s_logisimNet6),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus95[5:0]),
.dataB(s_logisimBus10[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_44
(.aEqualsB(s_logisimNet31),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus96[5:0]),
.dataB(s_logisimBus14[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_45
(.aEqualsB(s_logisimNet46),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus97[5:0]),
.dataB(s_logisimBus14[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_46
(.aEqualsB(s_logisimNet52),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus98[5:0]),
.dataB(s_logisimBus14[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_47
(.aEqualsB(s_logisimNet28),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus99[5:0]),
.dataB(s_logisimBus14[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_48
(.aEqualsB(s_logisimNet25),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus100[5:0]),
.dataB(s_logisimBus14[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_49
(.aEqualsB(s_logisimNet47),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus101[5:0]),
.dataB(s_logisimBus14[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_50
(.aEqualsB(s_logisimNet36),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus102[5:0]),
.dataB(s_logisimBus14[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_51
(.aEqualsB(s_logisimNet20),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus103[5:0]),
.dataB(s_logisimBus14[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_52
(.aEqualsB(s_logisimNet16),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus104[5:0]),
.dataB(s_logisimBus14[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_53
(.aEqualsB(s_logisimNet42),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus105[5:0]),
.dataB(s_logisimBus14[5:0]));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(1))
MEMORY_54
(.clock(s_logisimNet34),
.clockEnable(1'b1),
.d(s_logisimNet0),
.q(s_logisimNet7),
.reset(1'b0),
.tick(1'b1));
endmodule