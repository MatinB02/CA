/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
main
**
**
**
*****************************************************************************/
module
main(
InstDone,
Jen,
Jin,
Jout,
R1,
R10,
R11,
R12,
R13,
R14,
R15,
R16,
R17,
R18,
R19,
R2,
R20,
R21,
R22,
R23,
R24,
R25,
R26,
R27,
R28,
R29,
R3,
R30,
R31,
R4,
R5,
R6,
R7,
R8,
R9,
clk,
nop,
rst,
test
);
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
Jen;
input
[31:0]
Jin;
input
clk;
input
rst;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
InstDone;
output
[31:0]
Jout;
output
[31:0]
R1;
output
[31:0]
R10;
output
[31:0]
R11;
output
[31:0]
R12;
output
[31:0]
R13;
output
[31:0]
R14;
output
[31:0]
R15;
output
[31:0]
R16;
output
[31:0]
R17;
output
[31:0]
R18;
output
[31:0]
R19;
output
[31:0]
R2;
output
[31:0]
R20;
output
[31:0]
R21;
output
[31:0]
R22;
output
[31:0]
R23;
output
[31:0]
R24;
output
[31:0]
R25;
output
[31:0]
R26;
output
[31:0]
R27;
output
[31:0]
R28;
output
[31:0]
R29;
output
[31:0]
R3;
output
[31:0]
R30;
output
[31:0]
R31;
output
[31:0]
R4;
output
[31:0]
R5;
output
[31:0]
R6;
output
[31:0]
R7;
output
[31:0]
R8;
output
[31:0]
R9;
output
nop;
output
[31:0]
test;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
[31:0]
s_logisimBus0;
wire
[31:0]
s_logisimBus10;
wire
[4:0]
s_logisimBus11;
wire
[31:0]
s_logisimBus13;
wire
[15:0]
s_logisimBus14;
wire
[4:0]
s_logisimBus15;
wire
[8:0]
s_logisimBus16;
wire
[31:0]
s_logisimBus17;
wire
[5:0]
s_logisimBus18;
wire
[8:0]
s_logisimBus19;
wire
[31:0]
s_logisimBus20;
wire
[31:0]
s_logisimBus22;
wire
[31:0]
s_logisimBus23;
wire
[31:0]
s_logisimBus25;
wire
[4:0]
s_logisimBus27;
wire
[4:0]
s_logisimBus28;
wire
[31:0]
s_logisimBus29;
wire
[8:0]
s_logisimBus30;
wire
[4:0]
s_logisimBus31;
wire
[31:0]
s_logisimBus32;
wire
[31:0]
s_logisimBus33;
wire
[31:0]
s_logisimBus34;
wire
[31:0]
s_logisimBus38;
wire
[31:0]
s_logisimBus40;
wire
[31:0]
s_logisimBus41;
wire
[4:0]
s_logisimBus42;
wire
[8:0]
s_logisimBus43;
wire
[8:0]
s_logisimBus48;
wire
[31:0]
s_logisimBus49;
wire
[8:0]
s_logisimBus50;
wire
[4:0]
s_logisimBus54;
wire
[4:0]
s_logisimBus55;
wire
[31:0]
s_logisimBus56;
wire
[8:0]
s_logisimBus59;
wire
[3:0]
s_logisimBus6;
wire
[31:0]
s_logisimBus62;
wire
[31:0]
s_logisimBus67;
wire
[31:0]
s_logisimBus68;
wire
[31:0]
s_logisimBus69;
wire
[5:0]
s_logisimBus7;
wire
[31:0]
s_logisimBus70;
wire
[31:0]
s_logisimBus71;
wire
[31:0]
s_logisimBus72;
wire
[31:0]
s_logisimBus73;
wire
[31:0]
s_logisimBus74;
wire
[31:0]
s_logisimBus75;
wire
[31:0]
s_logisimBus76;
wire
[31:0]
s_logisimBus77;
wire
[31:0]
s_logisimBus78;
wire
[31:0]
s_logisimBus79;
wire
[31:0]
s_logisimBus80;
wire
[31:0]
s_logisimBus81;
wire
[31:0]
s_logisimBus82;
wire
[31:0]
s_logisimBus83;
wire
[31:0]
s_logisimBus84;
wire
[31:0]
s_logisimBus85;
wire
[31:0]
s_logisimBus86;
wire
[31:0]
s_logisimBus87;
wire
[31:0]
s_logisimBus88;
wire
[31:0]
s_logisimBus89;
wire
[4:0]
s_logisimBus9;
wire
[31:0]
s_logisimBus90;
wire
[31:0]
s_logisimBus91;
wire
[31:0]
s_logisimBus92;
wire
[31:0]
s_logisimBus93;
wire
[31:0]
s_logisimBus94;
wire
[31:0]
s_logisimBus95;
wire
[31:0]
s_logisimBus96;
wire
[31:0]
s_logisimBus97;
wire
[31:0]
s_logisimBus98;
wire
[31:0]
s_logisimBus99;
wire
s_logisimNet1;
wire
s_logisimNet12;
wire
s_logisimNet2;
wire
s_logisimNet21;
wire
s_logisimNet24;
wire
s_logisimNet26;
wire
s_logisimNet3;
wire
s_logisimNet35;
wire
s_logisimNet37;
wire
s_logisimNet39;
wire
s_logisimNet4;
wire
s_logisimNet44;
wire
s_logisimNet45;
wire
s_logisimNet46;
wire
s_logisimNet47;
wire
s_logisimNet5;
wire
s_logisimNet51;
wire
s_logisimNet52;
wire
s_logisimNet57;
wire
s_logisimNet60;
wire
s_logisimNet63;
wire
s_logisimNet64;
wire
s_logisimNet65;
wire
s_logisimNet66;
wire
s_logisimNet8;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
all
input
connections
are
defined
**
*******************************************************************************/
assign
s_logisimBus49[31:0]
=
Jin;
assign
s_logisimNet12
=
rst;
assign
s_logisimNet2
=
Jen;
assign
s_logisimNet47
=
clk;
/*******************************************************************************
**
Here
all
output
connections
are
defined
**
*******************************************************************************/
assign
InstDone
=
s_logisimNet26;
assign
Jout
=
s_logisimBus33[31:0];
assign
R1
=
s_logisimBus69[31:0];
assign
R10
=
s_logisimBus78[31:0];
assign
R11
=
s_logisimBus79[31:0];
assign
R12
=
s_logisimBus80[31:0];
assign
R13
=
s_logisimBus81[31:0];
assign
R14
=
s_logisimBus82[31:0];
assign
R15
=
s_logisimBus83[31:0];
assign
R16
=
s_logisimBus84[31:0];
assign
R17
=
s_logisimBus85[31:0];
assign
R18
=
s_logisimBus86[31:0];
assign
R19
=
s_logisimBus87[31:0];
assign
R2
=
s_logisimBus70[31:0];
assign
R20
=
s_logisimBus88[31:0];
assign
R21
=
s_logisimBus89[31:0];
assign
R22
=
s_logisimBus90[31:0];
assign
R23
=
s_logisimBus91[31:0];
assign
R24
=
s_logisimBus92[31:0];
assign
R25
=
s_logisimBus93[31:0];
assign
R26
=
s_logisimBus94[31:0];
assign
R27
=
s_logisimBus95[31:0];
assign
R28
=
s_logisimBus96[31:0];
assign
R29
=
s_logisimBus97[31:0];
assign
R3
=
s_logisimBus71[31:0];
assign
R30
=
s_logisimBus98[31:0];
assign
R31
=
s_logisimBus99[31:0];
assign
R4
=
s_logisimBus72[31:0];
assign
R5
=
s_logisimBus73[31:0];
assign
R6
=
s_logisimBus74[31:0];
assign
R7
=
s_logisimBus75[31:0];
assign
R8
=
s_logisimBus76[31:0];
assign
R9
=
s_logisimBus77[31:0];
assign
nop
=
s_logisimNet44;
assign
test
=
s_logisimBus32[31:0];
/*******************************************************************************
**
Here
all
in-lined
components
are
defined
**
*******************************************************************************/
assign
s_logisimBus13[0]
=
s_logisimBus11[0];
assign
s_logisimBus13[1]
=
s_logisimBus11[1];
assign
s_logisimBus13[2]
=
s_logisimBus11[2];
assign
s_logisimBus13[3]
=
s_logisimBus11[3];
assign
s_logisimBus13[4]
=
s_logisimBus11[4];
assign
s_logisimBus13[5]
=
1'b0;
assign
s_logisimBus13[6]
=
1'b0;
assign
s_logisimBus13[7]
=
1'b0;
assign
s_logisimBus13[8]
=
1'b0;
assign
s_logisimBus13[9]
=
1'b0;
assign
s_logisimBus13[10]
=
1'b0;
assign
s_logisimBus13[11]
=
1'b0;
assign
s_logisimBus13[12]
=
1'b0;
assign
s_logisimBus13[13]
=
1'b0;
assign
s_logisimBus13[14]
=
1'b0;
assign
s_logisimBus13[15]
=
1'b0;
assign
s_logisimBus13[16]
=
1'b0;
assign
s_logisimBus13[17]
=
1'b0;
assign
s_logisimBus13[18]
=
1'b0;
assign
s_logisimBus13[19]
=
1'b0;
assign
s_logisimBus13[20]
=
1'b0;
assign
s_logisimBus13[21]
=
1'b0;
assign
s_logisimBus13[22]
=
1'b0;
assign
s_logisimBus13[23]
=
1'b0;
assign
s_logisimBus13[24]
=
1'b0;
assign
s_logisimBus13[25]
=
1'b0;
assign
s_logisimBus13[26]
=
1'b0;
assign
s_logisimBus13[27]
=
1'b0;
assign
s_logisimBus13[28]
=
1'b0;
assign
s_logisimBus13[29]
=
1'b0;
assign
s_logisimBus13[30]
=
1'b0;
assign
s_logisimBus13[31]
=
1'b0;
assign
s_logisimBus59[8:0]
=
{1'b0,
8'h01};
assign
s_logisimBus54[4:0]
=
{1'b0,
4'h0};
assign
s_logisimBus55[4:0]
=
{1'b1,
4'hF};
assign
s_logisimBus56[0]
=
s_logisimBus50[0];
assign
s_logisimBus56[1]
=
s_logisimBus50[1];
assign
s_logisimBus56[2]
=
s_logisimBus50[2];
assign
s_logisimBus56[3]
=
s_logisimBus50[3];
assign
s_logisimBus56[4]
=
s_logisimBus50[4];
assign
s_logisimBus56[5]
=
s_logisimBus50[5];
assign
s_logisimBus56[6]
=
s_logisimBus50[6];
assign
s_logisimBus56[7]
=
s_logisimBus50[7];
assign
s_logisimBus56[8]
=
s_logisimBus50[8];
assign
s_logisimBus56[9]
=
s_logisimBus50[8];
assign
s_logisimBus56[10]
=
s_logisimBus50[8];
assign
s_logisimBus56[11]
=
s_logisimBus50[8];
assign
s_logisimBus56[12]
=
s_logisimBus50[8];
assign
s_logisimBus56[13]
=
s_logisimBus50[8];
assign
s_logisimBus56[14]
=
s_logisimBus50[8];
assign
s_logisimBus56[15]
=
s_logisimBus50[8];
assign
s_logisimBus56[16]
=
s_logisimBus50[8];
assign
s_logisimBus56[17]
=
s_logisimBus50[8];
assign
s_logisimBus56[18]
=
s_logisimBus50[8];
assign
s_logisimBus56[19]
=
s_logisimBus50[8];
assign
s_logisimBus56[20]
=
s_logisimBus50[8];
assign
s_logisimBus56[21]
=
s_logisimBus50[8];
assign
s_logisimBus56[22]
=
s_logisimBus50[8];
assign
s_logisimBus56[23]
=
s_logisimBus50[8];
assign
s_logisimBus56[24]
=
s_logisimBus50[8];
assign
s_logisimBus56[25]
=
s_logisimBus50[8];
assign
s_logisimBus56[26]
=
s_logisimBus50[8];
assign
s_logisimBus56[27]
=
s_logisimBus50[8];
assign
s_logisimBus56[28]
=
s_logisimBus50[8];
assign
s_logisimBus56[29]
=
s_logisimBus50[8];
assign
s_logisimBus56[30]
=
s_logisimBus50[8];
assign
s_logisimBus56[31]
=
s_logisimBus50[8];
assign
s_logisimBus34[0]
=
s_logisimBus14[0];
assign
s_logisimBus34[1]
=
s_logisimBus14[1];
assign
s_logisimBus34[2]
=
s_logisimBus14[2];
assign
s_logisimBus34[3]
=
s_logisimBus14[3];
assign
s_logisimBus34[4]
=
s_logisimBus14[4];
assign
s_logisimBus34[5]
=
s_logisimBus14[5];
assign
s_logisimBus34[6]
=
s_logisimBus14[6];
assign
s_logisimBus34[7]
=
s_logisimBus14[7];
assign
s_logisimBus34[8]
=
s_logisimBus14[8];
assign
s_logisimBus34[9]
=
s_logisimBus14[9];
assign
s_logisimBus34[10]
=
s_logisimBus14[10];
assign
s_logisimBus34[11]
=
s_logisimBus14[11];
assign
s_logisimBus34[12]
=
s_logisimBus14[12];
assign
s_logisimBus34[13]
=
s_logisimBus14[13];
assign
s_logisimBus34[14]
=
s_logisimBus14[14];
assign
s_logisimBus34[15]
=
s_logisimBus14[15];
assign
s_logisimBus34[16]
=
s_logisimBus14[15];
assign
s_logisimBus34[17]
=
s_logisimBus14[15];
assign
s_logisimBus34[18]
=
s_logisimBus14[15];
assign
s_logisimBus34[19]
=
s_logisimBus14[15];
assign
s_logisimBus34[20]
=
s_logisimBus14[15];
assign
s_logisimBus34[21]
=
s_logisimBus14[15];
assign
s_logisimBus34[22]
=
s_logisimBus14[15];
assign
s_logisimBus34[23]
=
s_logisimBus14[15];
assign
s_logisimBus34[24]
=
s_logisimBus14[15];
assign
s_logisimBus34[25]
=
s_logisimBus14[15];
assign
s_logisimBus34[26]
=
s_logisimBus14[15];
assign
s_logisimBus34[27]
=
s_logisimBus14[15];
assign
s_logisimBus34[28]
=
s_logisimBus14[15];
assign
s_logisimBus34[29]
=
s_logisimBus14[15];
assign
s_logisimBus34[30]
=
s_logisimBus14[15];
assign
s_logisimBus34[31]
=
s_logisimBus14[15];
/*******************************************************************************
**
Here
all
normal
components
are
defined
**
*******************************************************************************/
AND_GATE
#(.BubblesMask(2'b01))
GATES_1
(.input1(s_logisimNet35),
.input2(s_logisimNet64),
.result(s_logisimNet3));
OR_GATE
#(.BubblesMask(2'b00))
GATES_2
(.input1(s_logisimNet3),
.input2(s_logisimNet5),
.result(s_logisimNet24));
AND_GATE
#(.BubblesMask(2'b00))
GATES_3
(.input1(s_logisimNet35),
.input2(s_logisimNet66),
.result(s_logisimNet5));
OR_GATE
#(.BubblesMask(2'b00))
GATES_4
(.input1(s_logisimNet57),
.input2(s_logisimNet51),
.result(s_logisimNet52));
AND_GATE
#(.BubblesMask(2'b10))
GATES_5
(.input1(s_logisimNet47),
.input2(s_logisimNet44),
.result(s_logisimNet60));
Multiplexer_bus_2
#(.nrOfBits(32))
PLEXERS_6
(.enable(1'b1),
.muxIn_0(s_logisimBus17[31:0]),
.muxIn_1(s_logisimBus13[31:0]),
.muxOut(s_logisimBus41[31:0]),
.sel(s_logisimNet8));
Multiplexer_bus_2
#(.nrOfBits(32))
PLEXERS_7
(.enable(1'b1),
.muxIn_0(s_logisimBus67[31:0]),
.muxIn_1(s_logisimBus68[31:0]),
.muxOut(s_logisimBus10[31:0]),
.sel(s_logisimNet8));
Multiplexer_bus_2
#(.nrOfBits(9))
PLEXERS_8
(.enable(1'b1),
.muxIn_0(s_logisimBus50[8:0]),
.muxIn_1(s_logisimBus48[8:0]),
.muxOut(s_logisimBus43[8:0]),
.sel(s_logisimNet24));
Multiplexer_bus_2
#(.nrOfBits(9))
PLEXERS_9
(.enable(1'b1),
.muxIn_0(s_logisimBus43[8:0]),
.muxIn_1(s_logisimBus14[8:0]),
.muxOut(s_logisimBus19[8:0]),
.sel(s_logisimNet52));
Multiplexer_bus_2
#(.nrOfBits(9))
PLEXERS_10
(.enable(1'b1),
.muxIn_0(s_logisimBus19[8:0]),
.muxIn_1(s_logisimBus67[8:0]),
.muxOut(s_logisimBus30[8:0]),
.sel(s_logisimNet45));
Multiplexer_bus_2
#(.nrOfBits(5))
PLEXERS_11
(.enable(1'b1),
.muxIn_0(s_logisimBus31[4:0]),
.muxIn_1(s_logisimBus42[4:0]),
.muxOut(s_logisimBus27[4:0]),
.sel(s_logisimNet46));
Multiplexer_bus_2
#(.nrOfBits(32))
PLEXERS_12
(.enable(1'b1),
.muxIn_0(s_logisimBus40[31:0]),
.muxIn_1(s_logisimBus62[31:0]),
.muxOut(s_logisimBus0[31:0]),
.sel(s_logisimNet37));
Multiplexer_bus_2
#(.nrOfBits(5))
PLEXERS_13
(.enable(1'b1),
.muxIn_0(s_logisimBus54[4:0]),
.muxIn_1(s_logisimBus27[4:0]),
.muxOut(s_logisimBus15[4:0]),
.sel(s_logisimNet39));
Multiplexer_bus_2
#(.nrOfBits(32))
PLEXERS_14
(.enable(1'b1),
.muxIn_0(s_logisimBus0[31:0]),
.muxIn_1(s_logisimBus38[31:0]),
.muxOut(s_logisimBus22[31:0]),
.sel(s_logisimNet21));
Multiplexer_bus_2
#(.nrOfBits(5))
PLEXERS_15
(.enable(1'b1),
.muxIn_0(s_logisimBus15[4:0]),
.muxIn_1(s_logisimBus55[4:0]),
.muxOut(s_logisimBus9[4:0]),
.sel(s_logisimNet57));
Multiplexer_bus_2
#(.nrOfBits(32))
PLEXERS_16
(.enable(1'b1),
.muxIn_0(s_logisimBus22[31:0]),
.muxIn_1(s_logisimBus56[31:0]),
.muxOut(s_logisimBus20[31:0]),
.sel(s_logisimNet57));
Multiplexer_bus_2
#(.nrOfBits(32))
PLEXERS_17
(.enable(1'b1),
.muxIn_0(s_logisimBus68[31:0]),
.muxIn_1(s_logisimBus34[31:0]),
.muxOut(s_logisimBus17[31:0]),
.sel(s_logisimNet1));
Adder
#(.extendedBits(10),
.nrOfBits(9))
ARITH_18
(.carryIn(1'b0),
.carryOut(),
.dataA(s_logisimBus50[8:0]),
.dataB(s_logisimBus34[8:0]),
.result(s_logisimBus48[8:0]));
Adder
#(.extendedBits(10),
.nrOfBits(9))
ARITH_19
(.carryIn(1'b0),
.carryOut(),
.dataA(s_logisimBus16[8:0]),
.dataB(s_logisimBus59[8:0]),
.result(s_logisimBus50[8:0]));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(9))
pc
(.clock(s_logisimNet60),
.clockEnable(1'b1),
.d(s_logisimBus30[8:0]),
.q(s_logisimBus16[8:0]),
.reset(s_logisimNet12),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(32))
HI
(.clock(s_logisimNet60),
.clockEnable(s_logisimNet65),
.d(s_logisimBus29[31:0]),
.q(s_logisimBus38[31:0]),
.reset(1'b0),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(32))
LO
(.clock(s_logisimNet60),
.clockEnable(s_logisimNet65),
.d(s_logisimBus40[31:0]),
.q(s_logisimBus25[31:0]),
.reset(1'b0),
.tick(1'b1));
/*******************************************************************************
**
Here
all
sub-circuits
are
defined
**
*******************************************************************************/
jtag_ram512
Dmem
(.Addr(s_logisimBus40[8:0]),
.Din(s_logisimBus68[31:0]),
.Dout(s_logisimBus62[31:0]),
.Jen(s_logisimNet2),
.Jin(s_logisimBus23[31:0]),
.Jout(s_logisimBus33[31:0]),
.Wen(s_logisimNet63),
.clk(s_logisimNet60));
ALU
x3
(.InstDone(s_logisimNet26),
.a(s_logisimBus10[31:0]),
.aluop(s_logisimBus6[3:0]),
.b(s_logisimBus41[31:0]),
.clk(s_logisimNet47),
.res_high(s_logisimBus29[31:0]),
.res_low(s_logisimBus40[31:0]),
.zero(s_logisimNet35));
InstructionDecode
x1
(.Instruction(s_logisimBus32[31:0]),
.func(s_logisimBus18[5:0]),
.imm(s_logisimBus14[15:0]),
.opCode(s_logisimBus7[5:0]),
.rd(s_logisimBus42[4:0]),
.rs(s_logisimBus31[4:0]),
.rt(s_logisimBus28[4:0]),
.shmt(s_logisimBus11[4:0]));
ControlUnit
ControlUnit_1
(.ALUop(s_logisimBus6[3:0]),
.ALUsrc(s_logisimNet1),
.Rtype(),
.beq(s_logisimNet66),
.branch(s_logisimNet64),
.divv(s_logisimNet65),
.func(s_logisimBus18[5:0]),
.inst(s_logisimNet26),
.j(s_logisimNet51),
.jal(s_logisimNet57),
.jr(s_logisimNet45),
.main_clock(s_logisimNet47),
.memRead(),
.memToReg(s_logisimNet37),
.memWrite(s_logisimNet63),
.mohi(s_logisimNet21),
.mull(s_logisimNet4),
.nop(s_logisimNet44),
.opCode(s_logisimBus7[5:0]),
.regDst(s_logisimNet46),
.regWrite(s_logisimNet39),
.shmt(s_logisimNet8));
jtag_ram512
Imem
(.Addr(s_logisimBus16[8:0]),
.Din(32'd0),
.Dout(s_logisimBus32[31:0]),
.Jen(s_logisimNet2),
.Jin(s_logisimBus49[31:0]),
.Jout(s_logisimBus23[31:0]),
.Wen(1'b0),
.clk(s_logisimNet60));
regfile
x4
(.Aread0(s_logisimBus28[4:0]),
.Aread1(s_logisimBus31[4:0]),
.Awrite(s_logisimBus9[4:0]),
.Dread0(s_logisimBus67[31:0]),
.Dread1(s_logisimBus68[31:0]),
.Dwrite(s_logisimBus20[31:0]),
.R1(s_logisimBus69[31:0]),
.R10(s_logisimBus78[31:0]),
.R11(s_logisimBus79[31:0]),
.R12(s_logisimBus80[31:0]),
.R13(s_logisimBus81[31:0]),
.R14(s_logisimBus82[31:0]),
.R15(s_logisimBus83[31:0]),
.R16(s_logisimBus84[31:0]),
.R17(s_logisimBus85[31:0]),
.R18(s_logisimBus86[31:0]),
.R19(s_logisimBus87[31:0]),
.R2(s_logisimBus70[31:0]),
.R20(s_logisimBus88[31:0]),
.R21(s_logisimBus89[31:0]),
.R22(s_logisimBus90[31:0]),
.R23(s_logisimBus91[31:0]),
.R24(s_logisimBus92[31:0]),
.R25(s_logisimBus93[31:0]),
.R26(s_logisimBus94[31:0]),
.R27(s_logisimBus95[31:0]),
.R28(s_logisimBus96[31:0]),
.R29(s_logisimBus97[31:0]),
.R3(s_logisimBus71[31:0]),
.R30(s_logisimBus98[31:0]),
.R31(s_logisimBus99[31:0]),
.R4(s_logisimBus72[31:0]),
.R5(s_logisimBus73[31:0]),
.R6(s_logisimBus74[31:0]),
.R7(s_logisimBus75[31:0]),
.R8(s_logisimBus76[31:0]),
.R9(s_logisimBus77[31:0]),
.clk(s_logisimNet60),
.rst(s_logisimNet12));
endmodule