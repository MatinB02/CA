/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
ALU
**
**
**
*****************************************************************************/
module
ALU(
a,
aluop,
b,
res_high,
res_low
);
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
[31:0]
a;
input
[3:0]
aluop;
input
[31:0]
b;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
[31:0]
res_high;
output
[31:0]
res_low;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
[31:0]
s_logisimBus0;
wire
[31:0]
s_logisimBus1;
wire
[31:0]
s_logisimBus10;
wire
[31:0]
s_logisimBus12;
wire
[31:0]
s_logisimBus13;
wire
[31:0]
s_logisimBus14;
wire
[31:0]
s_logisimBus15;
wire
[31:0]
s_logisimBus16;
wire
[31:0]
s_logisimBus17;
wire
[31:0]
s_logisimBus18;
wire
[31:0]
s_logisimBus19;
wire
[31:0]
s_logisimBus2;
wire
[31:0]
s_logisimBus20;
wire
[3:0]
s_logisimBus21;
wire
[31:0]
s_logisimBus3;
wire
[31:0]
s_logisimBus4;
wire
[31:0]
s_logisimBus5;
wire
[31:0]
s_logisimBus6;
wire
[31:0]
s_logisimBus7;
wire
[3:0]
s_logisimBus8;
wire
[31:0]
s_logisimBus9;
wire
s_logisimNet11;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
all
input
connections
are
defined
**
*******************************************************************************/
assign
s_logisimBus3[31:0]
=
a;
assign
s_logisimBus6[31:0]
=
b;
assign
s_logisimBus8[3:0]
=
aluop;
/*******************************************************************************
**
Here
all
output
connections
are
defined
**
*******************************************************************************/
assign
res_high
=
s_logisimBus1[31:0];
assign
res_low
=
s_logisimBus15[31:0];
/*******************************************************************************
**
Here
all
in-lined
components
are
defined
**
*******************************************************************************/
assign
s_logisimBus21[3:0]
=
4'h1;
/*******************************************************************************
**
Here
all
normal
components
are
defined
**
*******************************************************************************/
Multiplexer_bus_16
#(.nrOfBits(32))
PLEXERS_1
(.enable(1'b1),
.muxIn_0(s_logisimBus0[31:0]),
.muxIn_1(s_logisimBus0[31:0]),
.muxIn_10(s_logisimBus9[31:0]),
.muxIn_11(s_logisimBus12[31:0]),
.muxIn_12(32'd0),
.muxIn_13(32'd0),
.muxIn_14(32'd0),
.muxIn_15(32'd0),
.muxIn_2(32'd0),
.muxIn_3(32'd0),
.muxIn_4(s_logisimBus4[31:0]),
.muxIn_5(s_logisimBus20[31:0]),
.muxIn_6(s_logisimBus2[31:0]),
.muxIn_7(32'd0),
.muxIn_8(32'd0),
.muxIn_9(s_logisimBus7[31:0]),
.muxOut(s_logisimBus1[31:0]),
.sel(s_logisimBus8[3:0]));
Multiplexer_bus_16
#(.nrOfBits(32))
PLEXERS_2
(.enable(1'b1),
.muxIn_0(s_logisimBus16[31:0]),
.muxIn_1(s_logisimBus16[31:0]),
.muxIn_10(s_logisimBus17[31:0]),
.muxIn_11(s_logisimBus18[31:0]),
.muxIn_12(s_logisimBus13[31:0]),
.muxIn_13(32'd0),
.muxIn_14(32'd0),
.muxIn_15(32'd0),
.muxIn_2(32'd0),
.muxIn_3(32'd0),
.muxIn_4(s_logisimBus5[31:0]),
.muxIn_5(s_logisimBus10[31:0]),
.muxIn_6(s_logisimBus19[31:0]),
.muxIn_7(32'd0),
.muxIn_8(32'd0),
.muxIn_9(s_logisimBus14[31:0]),
.muxOut(s_logisimBus15[31:0]),
.sel(s_logisimBus8[3:0]));
Comparator
#(.nrOfBits(4),
.twosComplement(0))
ARITH_3
(.aEqualsB(s_logisimNet11),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus8[3:0]),
.dataB(s_logisimBus21[3:0]));
Adder
#(.extendedBits(33),
.nrOfBits(32))
ARITH_4
(.carryIn(1'b0),
.carryOut(),
.dataA(s_logisimBus3[31:0]),
.dataB(s_logisimBus6[31:0]),
.result(s_logisimBus13[31:0]));
/*******************************************************************************
**
Here
all
sub-circuits
are
defined
**
*******************************************************************************/
ADDD
x1
(.S(s_logisimNet11),
.a(s_logisimBus3[31:0]),
.b(s_logisimBus6[31:0]),
.res_high(s_logisimBus0[31:0]),
.res_low(s_logisimBus16[31:0]));
ANDD
x2
(.a(s_logisimBus3[31:0]),
.b(s_logisimBus6[31:0]),
.res_high(s_logisimBus4[31:0]),
.res_low(s_logisimBus5[31:0]));
ORR
x3
(.a(s_logisimBus3[31:0]),
.b(s_logisimBus6[31:0]),
.res_high(s_logisimBus20[31:0]),
.res_low(s_logisimBus10[31:0]));
XORR
x4
(.a(s_logisimBus3[31:0]),
.b(s_logisimBus6[31:0]),
.res_high(s_logisimBus2[31:0]),
.res_low(s_logisimBus19[31:0]));
SLLL
x5
(.a(s_logisimBus3[31:0]),
.b(s_logisimBus6[31:0]),
.res_high(s_logisimBus7[31:0]),
.res_low(s_logisimBus14[31:0]));
SRLL
x6
(.a(s_logisimBus3[31:0]),
.b(s_logisimBus6[31:0]),
.res_high(s_logisimBus9[31:0]),
.res_low(s_logisimBus17[31:0]));
SRAA
x7
(.a(s_logisimBus3[31:0]),
.b(s_logisimBus6[31:0]),
.res_high(s_logisimBus12[31:0]),
.res_low(s_logisimBus18[31:0]));
endmodule