/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
MULL
**
**
**
*****************************************************************************/
module
MULL(
Done,
a,
b,
clk,
res_high,
res_low
);
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
[31:0]
a;
input
[31:0]
b;
input
clk;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
Done;
output
[31:0]
res_high;
output
[31:0]
res_low;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
[31:0]
s_logisimBus10;
wire
[31:0]
s_logisimBus11;
wire
[63:0]
s_logisimBus12;
wire
[31:0]
s_logisimBus13;
wire
[31:0]
s_logisimBus14;
wire
[7:0]
s_logisimBus15;
wire
[63:0]
s_logisimBus17;
wire
[7:0]
s_logisimBus18;
wire
[63:0]
s_logisimBus19;
wire
[63:0]
s_logisimBus2;
wire
[63:0]
s_logisimBus21;
wire
[63:0]
s_logisimBus22;
wire
[63:0]
s_logisimBus23;
wire
[63:0]
s_logisimBus28;
wire
[63:0]
s_logisimBus29;
wire
[63:0]
s_logisimBus3;
wire
[63:0]
s_logisimBus30;
wire
[31:0]
s_logisimBus31;
wire
[5:0]
s_logisimBus32;
wire
[31:0]
s_logisimBus33;
wire
[5:0]
s_logisimBus34;
wire
[7:0]
s_logisimBus37;
wire
[5:0]
s_logisimBus38;
wire
[63:0]
s_logisimBus4;
wire
[31:0]
s_logisimBus40;
wire
[63:0]
s_logisimBus5;
wire
[31:0]
s_logisimBus7;
wire
[63:0]
s_logisimBus8;
wire
s_logisimNet0;
wire
s_logisimNet1;
wire
s_logisimNet16;
wire
s_logisimNet20;
wire
s_logisimNet25;
wire
s_logisimNet26;
wire
s_logisimNet27;
wire
s_logisimNet36;
wire
s_logisimNet39;
wire
s_logisimNet6;
wire
s_logisimNet9;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
all
input
connections
are
defined
**
*******************************************************************************/
assign
s_logisimBus10[31:0]
=
b;
assign
s_logisimBus11[31:0]
=
a;
assign
s_logisimNet9
=
clk;
/*******************************************************************************
**
Here
all
output
connections
are
defined
**
*******************************************************************************/
assign
Done
=
s_logisimNet16;
assign
res_high
=
s_logisimBus3[63:32];
assign
res_low
=
s_logisimBus3[31:0];
/*******************************************************************************
**
Here
all
in-lined
components
are
defined
**
*******************************************************************************/
assign
s_logisimBus5[63:0]
=
64'h0000000000000000;
assign
s_logisimBus34[5:0]
=
{2'b00,
4'h1};
assign
s_logisimBus18[7:0]
=
8'h10;
assign
s_logisimBus40[31:0]
=
32'h00000002;
assign
s_logisimBus37[7:0]
=
8'h01;
assign
s_logisimBus30[0]
=
s_logisimBus11[0];
assign
s_logisimBus30[1]
=
s_logisimBus11[1];
assign
s_logisimBus30[2]
=
s_logisimBus11[2];
assign
s_logisimBus30[3]
=
s_logisimBus11[3];
assign
s_logisimBus30[4]
=
s_logisimBus11[4];
assign
s_logisimBus30[5]
=
s_logisimBus11[5];
assign
s_logisimBus30[6]
=
s_logisimBus11[6];
assign
s_logisimBus30[7]
=
s_logisimBus11[7];
assign
s_logisimBus30[8]
=
s_logisimBus11[8];
assign
s_logisimBus30[9]
=
s_logisimBus11[9];
assign
s_logisimBus30[10]
=
s_logisimBus11[10];
assign
s_logisimBus30[11]
=
s_logisimBus11[11];
assign
s_logisimBus30[12]
=
s_logisimBus11[12];
assign
s_logisimBus30[13]
=
s_logisimBus11[13];
assign
s_logisimBus30[14]
=
s_logisimBus11[14];
assign
s_logisimBus30[15]
=
s_logisimBus11[15];
assign
s_logisimBus30[16]
=
s_logisimBus11[16];
assign
s_logisimBus30[17]
=
s_logisimBus11[17];
assign
s_logisimBus30[18]
=
s_logisimBus11[18];
assign
s_logisimBus30[19]
=
s_logisimBus11[19];
assign
s_logisimBus30[20]
=
s_logisimBus11[20];
assign
s_logisimBus30[21]
=
s_logisimBus11[21];
assign
s_logisimBus30[22]
=
s_logisimBus11[22];
assign
s_logisimBus30[23]
=
s_logisimBus11[23];
assign
s_logisimBus30[24]
=
s_logisimBus11[24];
assign
s_logisimBus30[25]
=
s_logisimBus11[25];
assign
s_logisimBus30[26]
=
s_logisimBus11[26];
assign
s_logisimBus30[27]
=
s_logisimBus11[27];
assign
s_logisimBus30[28]
=
s_logisimBus11[28];
assign
s_logisimBus30[29]
=
s_logisimBus11[29];
assign
s_logisimBus30[30]
=
s_logisimBus11[30];
assign
s_logisimBus30[31]
=
s_logisimBus11[31];
assign
s_logisimBus30[32]
=
1'b0;
assign
s_logisimBus30[33]
=
1'b0;
assign
s_logisimBus30[34]
=
1'b0;
assign
s_logisimBus30[35]
=
1'b0;
assign
s_logisimBus30[36]
=
1'b0;
assign
s_logisimBus30[37]
=
1'b0;
assign
s_logisimBus30[38]
=
1'b0;
assign
s_logisimBus30[39]
=
1'b0;
assign
s_logisimBus30[40]
=
1'b0;
assign
s_logisimBus30[41]
=
1'b0;
assign
s_logisimBus30[42]
=
1'b0;
assign
s_logisimBus30[43]
=
1'b0;
assign
s_logisimBus30[44]
=
1'b0;
assign
s_logisimBus30[45]
=
1'b0;
assign
s_logisimBus30[46]
=
1'b0;
assign
s_logisimBus30[47]
=
1'b0;
assign
s_logisimBus30[48]
=
1'b0;
assign
s_logisimBus30[49]
=
1'b0;
assign
s_logisimBus30[50]
=
1'b0;
assign
s_logisimBus30[51]
=
1'b0;
assign
s_logisimBus30[52]
=
1'b0;
assign
s_logisimBus30[53]
=
1'b0;
assign
s_logisimBus30[54]
=
1'b0;
assign
s_logisimBus30[55]
=
1'b0;
assign
s_logisimBus30[56]
=
1'b0;
assign
s_logisimBus30[57]
=
1'b0;
assign
s_logisimBus30[58]
=
1'b0;
assign
s_logisimBus30[59]
=
1'b0;
assign
s_logisimBus30[60]
=
1'b0;
assign
s_logisimBus30[61]
=
1'b0;
assign
s_logisimBus30[62]
=
1'b0;
assign
s_logisimBus30[63]
=
1'b0;
assign
s_logisimBus32[5:0]
=
{2'b00,
4'h1};
assign
s_logisimBus38[5:0]
=
{2'b00,
4'h1};
assign
s_logisimNet36
=
~s_logisimNet1;
/*******************************************************************************
**
Here
all
normal
components
are
defined
**
*******************************************************************************/
NAND_GATE
#(.BubblesMask(2'b00))
GATES_1
(.input1(s_logisimNet27),
.input2(s_logisimNet26),
.result(s_logisimNet6));
OR_GATE
#(.BubblesMask(2'b00))
GATES_2
(.input1(s_logisimNet16),
.input2(s_logisimNet36),
.result(s_logisimNet39));
Multiplexer_bus_2
#(.nrOfBits(64))
PLEXERS_3
(.enable(1'b1),
.muxIn_0(s_logisimBus5[63:0]),
.muxIn_1(s_logisimBus12[63:0]),
.muxOut(s_logisimBus4[63:0]),
.sel(s_logisimBus14[0]));
Multiplexer_bus_2
#(.nrOfBits(64))
PLEXERS_4
(.enable(1'b1),
.muxIn_0(s_logisimBus5[63:0]),
.muxIn_1(s_logisimBus29[63:0]),
.muxOut(s_logisimBus22[63:0]),
.sel(s_logisimBus14[1]));
Multiplexer_bus_2
#(.nrOfBits(32))
PLEXERS_5
(.enable(1'b1),
.muxIn_0(s_logisimBus13[31:0]),
.muxIn_1(s_logisimBus10[31:0]),
.muxOut(s_logisimBus31[31:0]),
.sel(s_logisimNet6));
Multiplexer_bus_2
#(.nrOfBits(64))
PLEXERS_6
(.enable(1'b1),
.muxIn_0(s_logisimBus23[63:0]),
.muxIn_1(s_logisimBus30[63:0]),
.muxOut(s_logisimBus2[63:0]),
.sel(s_logisimNet6));
Shifter_64_bit
#(.shifterMode(0))
ARITH_7
(.dataA(s_logisimBus28[63:0]),
.result(s_logisimBus8[63:0]),
.shiftAmount(s_logisimBus34[5:0]));
Adder
#(.extendedBits(65),
.nrOfBits(64))
ARITH_8
(.carryIn(1'b0),
.carryOut(),
.dataA(s_logisimBus17[63:0]),
.dataB(s_logisimBus8[63:0]),
.result(s_logisimBus19[63:0]));
Comparator
#(.nrOfBits(32),
.twosComplement(1))
ARITH_9
(.aEqualsB(s_logisimNet27),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus33[31:0]),
.dataB(s_logisimBus10[31:0]));
Comparator
#(.nrOfBits(32),
.twosComplement(1))
ARITH_10
(.aEqualsB(s_logisimNet26),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus7[31:0]),
.dataB(s_logisimBus11[31:0]));
Comparator
#(.nrOfBits(8),
.twosComplement(1))
ARITH_11
(.aEqualsB(),
.aGreaterThanB(),
.aLessThanB(s_logisimNet1),
.dataA(s_logisimBus37[7:0]),
.dataB(s_logisimBus15[7:0]));
Shifter_64_bit
#(.shifterMode(0))
ARITH_12
(.dataA(s_logisimBus2[63:0]),
.result(s_logisimBus21[63:0]),
.shiftAmount(s_logisimBus32[5:0]));
Shifter_64_bit
#(.shifterMode(0))
ARITH_13
(.dataA(s_logisimBus29[63:0]),
.result(s_logisimBus23[63:0]),
.shiftAmount(s_logisimBus38[5:0]));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(32))
MEMORY_14
(.clock(s_logisimNet9),
.clockEnable(1'b1),
.d(s_logisimBus10[31:0]),
.q(s_logisimBus33[31:0]),
.reset(1'b0),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(32))
MEMORY_15
(.clock(s_logisimNet9),
.clockEnable(1'b1),
.d(s_logisimBus11[31:0]),
.q(s_logisimBus7[31:0]),
.reset(1'b0),
.tick(1'b1));
LogisimCounter
#(.invertClock(0),
.maxVal(8'hFF),
.mode(0),
.width(8))
MEMORY_16
(.clear(1'b0),
.clock(s_logisimNet9),
.compareOut(),
.countValue(s_logisimBus15[7:0]),
.enable(1'b1),
.load(s_logisimNet6),
.loadData(s_logisimBus18[7:0]),
.tick(1'b1),
.upNotDown(1'b0));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(32))
bb
(.clock(s_logisimNet9),
.clockEnable(s_logisimNet0),
.d(s_logisimBus31[31:0]),
.q(s_logisimBus14[31:0]),
.reset(1'b0),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(64))
aa
(.clock(s_logisimNet9),
.clockEnable(s_logisimNet0),
.d(s_logisimBus2[63:0]),
.q(s_logisimBus12[63:0]),
.reset(1'b0),
.tick(1'b1));
D_FLIPFLOP
#(.invertClockEnable(0))
MEMORY_19
(.clock(s_logisimNet9),
.d(s_logisimNet39),
.preset(1'b0),
.q(s_logisimNet16),
.qBar(s_logisimNet0),
.reset(s_logisimNet6),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(64))
aa1
(.clock(s_logisimNet9),
.clockEnable(s_logisimNet0),
.d(s_logisimBus21[63:0]),
.q(s_logisimBus29[63:0]),
.reset(1'b0),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(64))
P
(.clock(s_logisimNet9),
.clockEnable(s_logisimNet0),
.d(s_logisimBus19[63:0]),
.q(s_logisimBus3[63:0]),
.reset(s_logisimNet6),
.tick(1'b1));
/*******************************************************************************
**
Here
all
sub-circuits
are
defined
**
*******************************************************************************/
FAA
FAA_1
(.a(s_logisimBus4[63:0]),
.b(s_logisimBus22[63:0]),
.c(s_logisimBus3[63:0]),
.cout(s_logisimBus28[63:0]),
.s(s_logisimBus17[63:0]));
SRLL
SRLL_1
(.a(s_logisimBus14[31:0]),
.b(s_logisimBus40[31:0]),
.res_high(),
.res_low(s_logisimBus13[31:0]));
endmodule