/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
ControlUnit
**
**
**
*****************************************************************************/
module
ControlUnit(
ALUop,
ALUsrc,
addi_lw,
beq,
branchN,
clock,
func,
j,
jal,
jr,
link,
memToReg,
memWrite,
opCode,
regDst,
regWrite,
rst,
shift
);
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
clock;
input
[5:0]
func;
input
[5:0]
opCode;
input
rst;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
[3:0]
ALUop;
output
ALUsrc;
output
addi_lw;
output
beq;
output
branchN;
output
j;
output
jal;
output
jr;
output
link;
output
memToReg;
output
memWrite;
output
regDst;
output
regWrite;
output
shift;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
[3:0]
s_logisimBus14;
wire
[5:0]
s_logisimBus2;
wire
[5:0]
s_logisimBus3;
wire
[5:0]
s_logisimBus4;
wire
[5:0]
s_logisimBus5;
wire
[5:0]
s_logisimBus6;
wire
[5:0]
s_logisimBus7;
wire
[5:0]
s_logisimBus8;
wire
[5:0]
s_logisimBus9;
wire
s_logisimNet0;
wire
s_logisimNet1;
wire
s_logisimNet10;
wire
s_logisimNet11;
wire
s_logisimNet12;
wire
s_logisimNet13;
wire
s_logisimNet15;
wire
s_logisimNet16;
wire
s_logisimNet17;
wire
s_logisimNet18;
wire
s_logisimNet19;
wire
s_logisimNet20;
wire
s_logisimNet21;
wire
s_logisimNet22;
wire
s_logisimNet23;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
all
input
connections
are
defined
**
*******************************************************************************/
assign
s_logisimBus3[5:0]
=
func;
assign
s_logisimBus7[5:0]
=
opCode;
assign
s_logisimNet0
=
clock;
assign
s_logisimNet1
=
rst;
/*******************************************************************************
**
Here
all
output
connections
are
defined
**
*******************************************************************************/
assign
ALUop
=
s_logisimBus14[3:0];
assign
ALUsrc
=
s_logisimNet17;
assign
addi_lw
=
s_logisimNet23;
assign
beq
=
s_logisimNet22;
assign
branchN
=
s_logisimNet19;
assign
j
=
s_logisimNet16;
assign
jal
=
s_logisimNet21;
assign
jr
=
s_logisimNet20;
assign
link
=
s_logisimNet13;
assign
memToReg
=
s_logisimNet12;
assign
memWrite
=
s_logisimNet10;
assign
regDst
=
s_logisimNet15;
assign
regWrite
=
s_logisimNet11;
assign
shift
=
s_logisimNet18;
/*******************************************************************************
**
Here
all
normal
components
are
defined
**
*******************************************************************************/
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(6))
MEMORY_1
(.clock(s_logisimNet0),
.clockEnable(1'b1),
.d(s_logisimBus2[5:0]),
.q(s_logisimBus5[5:0]),
.reset(s_logisimNet1),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(6))
MEMORY_2
(.clock(s_logisimNet0),
.clockEnable(1'b1),
.d(s_logisimBus9[5:0]),
.q(s_logisimBus8[5:0]),
.reset(s_logisimNet1),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(6))
MEMORY_3
(.clock(s_logisimNet0),
.clockEnable(1'b1),
.d(s_logisimBus7[5:0]),
.q(s_logisimBus6[5:0]),
.reset(s_logisimNet1),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(6))
MEMORY_4
(.clock(s_logisimNet0),
.clockEnable(1'b1),
.d(s_logisimBus3[5:0]),
.q(s_logisimBus4[5:0]),
.reset(s_logisimNet1),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(6))
MEMORY_5
(.clock(s_logisimNet0),
.clockEnable(1'b1),
.d(s_logisimBus6[5:0]),
.q(s_logisimBus2[5:0]),
.reset(s_logisimNet1),
.tick(1'b1));
REGISTER_FLIP_FLOP
#(.invertClock(0),
.nrOfBits(6))
MEMORY_6
(.clock(s_logisimNet0),
.clockEnable(1'b1),
.d(s_logisimBus4[5:0]),
.q(s_logisimBus9[5:0]),
.reset(s_logisimNet1),
.tick(1'b1));
/*******************************************************************************
**
Here
all
sub-circuits
are
defined
**
*******************************************************************************/
CU4
CU4_1
(.memWrite(s_logisimNet10),
.opCode(s_logisimBus2[5:0]));
CU5
CU5_1
(.func(s_logisimBus8[5:0]),
.link(s_logisimNet13),
.memToReg(s_logisimNet12),
.opCode(s_logisimBus5[5:0]),
.regWrite(s_logisimNet11));
CU3
CU3_1
(.ALUop(s_logisimBus14[3:0]),
.ALUsrc(s_logisimNet17),
.addi_lw(s_logisimNet23),
.beq(s_logisimNet22),
.branchN(s_logisimNet19),
.func(s_logisimBus4[5:0]),
.j(s_logisimNet16),
.jal(s_logisimNet21),
.jr(s_logisimNet20),
.opCode(s_logisimBus6[5:0]),
.regDst(s_logisimNet15),
.shift(s_logisimNet18));
endmodule