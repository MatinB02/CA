/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
FP_ALU
**
**
**
*****************************************************************************/
module
FP_ALU(
Done,
a,
aluop,
b,
clk,
fsin,
res
);
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
[31:0]
a;
input
[2:0]
aluop;
input
[31:0]
b;
input
clk;
input
fsin;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
Done;
output
[31:0]
res;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
[31:0]
s_logisimBus0;
wire
[31:0]
s_logisimBus1;
wire
[31:0]
s_logisimBus13;
wire
[31:0]
s_logisimBus15;
wire
[31:0]
s_logisimBus2;
wire
[2:0]
s_logisimBus3;
wire
[31:0]
s_logisimBus5;
wire
[31:0]
s_logisimBus6;
wire
[31:0]
s_logisimBus7;
wire
[31:0]
s_logisimBus8;
wire
[2:0]
s_logisimBus9;
wire
s_logisimNet10;
wire
s_logisimNet11;
wire
s_logisimNet12;
wire
s_logisimNet14;
wire
s_logisimNet16;
wire
s_logisimNet4;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
all
input
connections
are
defined
**
*******************************************************************************/
assign
s_logisimBus0[31:0]
=
b;
assign
s_logisimBus3[2:0]
=
aluop;
assign
s_logisimBus7[31:0]
=
a;
assign
s_logisimNet11
=
clk;
assign
s_logisimNet16
=
fsin;
/*******************************************************************************
**
Here
all
output
connections
are
defined
**
*******************************************************************************/
assign
Done
=
s_logisimNet10;
assign
res
=
s_logisimBus13[31:0];
/*******************************************************************************
**
Here
all
in-lined
components
are
defined
**
*******************************************************************************/
assign
s_logisimBus9[2:0]
=
3'b101;
assign
s_logisimNet14
=
1'b1;
/*******************************************************************************
**
Here
all
normal
components
are
defined
**
*******************************************************************************/
Multiplexer_bus_8
#(.nrOfBits(32))
PLEXERS_1
(.enable(1'b1),
.muxIn_0(s_logisimBus2[31:0]),
.muxIn_1(s_logisimBus1[31:0]),
.muxIn_2(s_logisimBus8[31:0]),
.muxIn_3(s_logisimBus5[31:0]),
.muxIn_4(s_logisimBus15[31:0]),
.muxIn_5(s_logisimBus6[31:0]),
.muxIn_6(32'd0),
.muxIn_7(32'd0),
.muxOut(s_logisimBus13[31:0]),
.sel(s_logisimBus3[2:0]));
Multiplexer_2
PLEXERS_2
(.enable(1'b1),
.muxIn_0(s_logisimNet14),
.muxIn_1(s_logisimNet4),
.muxOut(s_logisimNet10),
.sel(s_logisimNet12));
Comparator
#(.nrOfBits(3),
.twosComplement(0))
ARITH_3
(.aEqualsB(s_logisimNet12),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus3[2:0]),
.dataB(s_logisimBus9[2:0]));
/*******************************************************************************
**
Here
all
sub-circuits
are
defined
**
*******************************************************************************/
fadd
faddH
(.INFINITY_PIN(),
.NAN_PIN(),
.a(s_logisimBus7[31:0]),
.b(s_logisimBus0[31:0]),
.res(s_logisimBus2[31:0]));
fsub
fsubH
(.INFINITY_PIN(),
.NAN_PIN(),
.a(s_logisimBus7[31:0]),
.b(s_logisimBus0[31:0]),
.res(s_logisimBus1[31:0]));
fmult
fmultH
(.a(s_logisimBus0[31:0]),
.b(s_logisimBus7[31:0]),
.res(s_logisimBus8[31:0]));
fabs
fabsH
(.a(s_logisimBus7[31:0]),
.res(s_logisimBus5[31:0]));
fslt
fsltH
(.INFINITY_PIN(),
.NAN_PIN(),
.a(s_logisimBus7[31:0]),
.b(s_logisimBus0[31:0]),
.res(s_logisimBus15[31:0]));
fsinn
fsinH
(.a(s_logisimBus7[31:0]),
.b(s_logisimBus0[31:0]),
.clk(s_logisimNet11),
.done(s_logisimNet4),
.fsin(s_logisimNet16),
.res(s_logisimBus6[31:0]));
endmodule