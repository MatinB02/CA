/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
CU3
**
**
**
*****************************************************************************/
module
CU3(
ALUop,
ALUsrc,
addi_lw,
beq,
branchN,
func,
j,
jal,
jr,
opCode,
regDst,
shift
);
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
[5:0]
func;
input
[5:0]
opCode;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
[3:0]
ALUop;
output
ALUsrc;
output
addi_lw;
output
beq;
output
branchN;
output
j;
output
jal;
output
jr;
output
regDst;
output
shift;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
[3:0]
s_logisimBus10;
wire
[3:0]
s_logisimBus11;
wire
[3:0]
s_logisimBus13;
wire
[3:0]
s_logisimBus14;
wire
[5:0]
s_logisimBus15;
wire
[3:0]
s_logisimBus16;
wire
[3:0]
s_logisimBus18;
wire
[3:0]
s_logisimBus23;
wire
[3:0]
s_logisimBus24;
wire
[3:0]
s_logisimBus25;
wire
[3:0]
s_logisimBus26;
wire
[3:0]
s_logisimBus30;
wire
[3:0]
s_logisimBus33;
wire
[3:0]
s_logisimBus34;
wire
[3:0]
s_logisimBus35;
wire
[3:0]
s_logisimBus37;
wire
[3:0]
s_logisimBus38;
wire
[3:0]
s_logisimBus39;
wire
[3:0]
s_logisimBus40;
wire
[3:0]
s_logisimBus49;
wire
[3:0]
s_logisimBus50;
wire
[3:0]
s_logisimBus51;
wire
[3:0]
s_logisimBus52;
wire
[3:0]
s_logisimBus53;
wire
[3:0]
s_logisimBus54;
wire
[3:0]
s_logisimBus55;
wire
[3:0]
s_logisimBus56;
wire
[3:0]
s_logisimBus57;
wire
[3:0]
s_logisimBus58;
wire
[3:0]
s_logisimBus59;
wire
[3:0]
s_logisimBus60;
wire
[3:0]
s_logisimBus61;
wire
[3:0]
s_logisimBus62;
wire
[3:0]
s_logisimBus63;
wire
[3:0]
s_logisimBus64;
wire
[3:0]
s_logisimBus65;
wire
[3:0]
s_logisimBus66;
wire
[3:0]
s_logisimBus67;
wire
[3:0]
s_logisimBus68;
wire
[3:0]
s_logisimBus69;
wire
[3:0]
s_logisimBus7;
wire
[5:0]
s_logisimBus70;
wire
[5:0]
s_logisimBus72;
wire
[5:0]
s_logisimBus73;
wire
[5:0]
s_logisimBus74;
wire
[5:0]
s_logisimBus75;
wire
[5:0]
s_logisimBus76;
wire
[5:0]
s_logisimBus77;
wire
[5:0]
s_logisimBus78;
wire
[5:0]
s_logisimBus79;
wire
[3:0]
s_logisimBus8;
wire
[5:0]
s_logisimBus80;
wire
[5:0]
s_logisimBus81;
wire
[5:0]
s_logisimBus82;
wire
[5:0]
s_logisimBus83;
wire
[5:0]
s_logisimBus84;
wire
[5:0]
s_logisimBus85;
wire
[5:0]
s_logisimBus86;
wire
[5:0]
s_logisimBus87;
wire
[5:0]
s_logisimBus88;
wire
[5:0]
s_logisimBus89;
wire
[5:0]
s_logisimBus9;
wire
[5:0]
s_logisimBus90;
wire
[5:0]
s_logisimBus91;
wire
[5:0]
s_logisimBus92;
wire
[5:0]
s_logisimBus93;
wire
[5:0]
s_logisimBus94;
wire
s_logisimNet0;
wire
s_logisimNet1;
wire
s_logisimNet12;
wire
s_logisimNet17;
wire
s_logisimNet19;
wire
s_logisimNet2;
wire
s_logisimNet20;
wire
s_logisimNet21;
wire
s_logisimNet22;
wire
s_logisimNet27;
wire
s_logisimNet28;
wire
s_logisimNet29;
wire
s_logisimNet3;
wire
s_logisimNet31;
wire
s_logisimNet32;
wire
s_logisimNet36;
wire
s_logisimNet4;
wire
s_logisimNet41;
wire
s_logisimNet42;
wire
s_logisimNet43;
wire
s_logisimNet44;
wire
s_logisimNet45;
wire
s_logisimNet46;
wire
s_logisimNet47;
wire
s_logisimNet48;
wire
s_logisimNet5;
wire
s_logisimNet6;
wire
s_logisimNet71;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
all
input
connections
are
defined
**
*******************************************************************************/
assign
s_logisimBus15[5:0]
=
func;
assign
s_logisimBus9[5:0]
=
opCode;
/*******************************************************************************
**
Here
all
output
connections
are
defined
**
*******************************************************************************/
assign
ALUop
=
s_logisimBus30[3:0];
assign
ALUsrc
=
s_logisimNet47;
assign
addi_lw
=
s_logisimNet17;
assign
beq
=
s_logisimNet44;
assign
branchN
=
s_logisimNet43;
assign
j
=
s_logisimNet6;
assign
jal
=
s_logisimNet22;
assign
jr
=
s_logisimNet19;
assign
regDst
=
s_logisimNet48;
assign
shift
=
s_logisimNet41;
/*******************************************************************************
**
Here
all
in-lined
components
are
defined
**
*******************************************************************************/
assign
s_logisimBus70[5:0]
=
{2'b10,
4'h0};
assign
s_logisimBus72[5:0]
=
{2'b10,
4'h2};
assign
s_logisimBus73[5:0]
=
{2'b10,
4'h4};
assign
s_logisimBus74[5:0]
=
{2'b10,
4'h5};
assign
s_logisimBus75[5:0]
=
{2'b10,
4'h6};
assign
s_logisimBus76[5:0]
=
{2'b00,
4'h4};
assign
s_logisimBus77[5:0]
=
{2'b00,
4'h6};
assign
s_logisimBus78[5:0]
=
{2'b00,
4'h7};
assign
s_logisimBus79[5:0]
=
{2'b01,
4'hA};
assign
s_logisimBus80[5:0]
=
{2'b01,
4'h0};
assign
s_logisimBus81[5:0]
=
{2'b00,
4'h0};
assign
s_logisimBus82[5:0]
=
{2'b00,
4'h8};
assign
s_logisimBus83[5:0]
=
{2'b01,
4'h2};
assign
s_logisimBus84[5:0]
=
{2'b00,
4'h2};
assign
s_logisimBus49[3:0]
=
4'h0;
assign
s_logisimBus50[3:0]
=
4'h1;
assign
s_logisimBus51[3:0]
=
4'h4;
assign
s_logisimBus52[3:0]
=
4'h5;
assign
s_logisimBus53[3:0]
=
4'h6;
assign
s_logisimBus85[5:0]
=
{2'b00,
4'h0};
assign
s_logisimBus86[5:0]
=
{2'b00,
4'h8};
assign
s_logisimBus87[5:0]
=
{2'b10,
4'hB};
assign
s_logisimBus88[5:0]
=
{2'b10,
4'h3};
assign
s_logisimBus89[5:0]
=
{2'b00,
4'h5};
assign
s_logisimBus90[5:0]
=
{2'b00,
4'hA};
assign
s_logisimBus91[5:0]
=
{2'b00,
4'h2};
assign
s_logisimBus92[5:0]
=
{2'b00,
4'h3};
assign
s_logisimBus93[5:0]
=
{2'b00,
4'h4};
assign
s_logisimBus94[5:0]
=
{2'b01,
4'hC};
assign
s_logisimBus54[3:0]
=
4'h9;
assign
s_logisimBus55[3:0]
=
4'hA;
assign
s_logisimBus56[3:0]
=
4'hB;
assign
s_logisimBus57[3:0]
=
4'h3;
assign
s_logisimBus58[3:0]
=
4'hF;
assign
s_logisimBus59[3:0]
=
4'h9;
assign
s_logisimBus60[3:0]
=
4'hF;
assign
s_logisimBus61[3:0]
=
4'hF;
assign
s_logisimBus62[3:0]
=
4'hC;
assign
s_logisimBus63[3:0]
=
4'h0;
assign
s_logisimBus64[3:0]
=
4'h0;
assign
s_logisimBus65[3:0]
=
4'h7;
assign
s_logisimBus66[3:0]
=
4'h2;
assign
s_logisimBus67[3:0]
=
4'hF;
assign
s_logisimBus68[3:0]
=
4'h1;
assign
s_logisimBus69[3:0]
=
4'h8;
/*******************************************************************************
**
Here
all
normal
components
are
defined
**
*******************************************************************************/
OR_GATE
#(.BubblesMask(2'b00))
GATES_1
(.input1(s_logisimNet27),
.input2(s_logisimNet29),
.result(s_logisimNet17));
AND_GATE
#(.BubblesMask(2'b00))
GATES_2
(.input1(s_logisimNet3),
.input2(s_logisimNet46),
.result(s_logisimNet45));
OR_GATE_5_INPUTS
#(.BubblesMask({1'b0,
4'h0}))
GATES_3
(.input1(s_logisimNet27),
.input2(s_logisimNet42),
.input3(s_logisimNet29),
.input4(s_logisimNet43),
.input5(s_logisimNet36),
.result(s_logisimNet47));
OR_GATE
#(.BubblesMask(2'b00))
GATES_4
(.input1(s_logisimNet45),
.input2(s_logisimNet31),
.result(s_logisimNet48));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_5
(.enable(1'b1),
.muxIn_0(s_logisimBus49[3:0]),
.muxIn_1(s_logisimBus50[3:0]),
.muxOut(s_logisimBus37[3:0]),
.sel(s_logisimNet4));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_6
(.enable(1'b1),
.muxIn_0(s_logisimBus37[3:0]),
.muxIn_1(s_logisimBus51[3:0]),
.muxOut(s_logisimBus23[3:0]),
.sel(s_logisimNet5));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_7
(.enable(1'b1),
.muxIn_0(s_logisimBus23[3:0]),
.muxIn_1(s_logisimBus52[3:0]),
.muxOut(s_logisimBus14[3:0]),
.sel(s_logisimNet12));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_8
(.enable(1'b1),
.muxIn_0(s_logisimBus14[3:0]),
.muxIn_1(s_logisimBus53[3:0]),
.muxOut(s_logisimBus13[3:0]),
.sel(s_logisimNet21));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_9
(.enable(1'b1),
.muxIn_0(s_logisimBus13[3:0]),
.muxIn_1(s_logisimBus54[3:0]),
.muxOut(s_logisimBus40[3:0]),
.sel(s_logisimNet2));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_10
(.enable(1'b1),
.muxIn_0(s_logisimBus40[3:0]),
.muxIn_1(s_logisimBus55[3:0]),
.muxOut(s_logisimBus26[3:0]),
.sel(s_logisimNet32));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_11
(.enable(1'b1),
.muxIn_0(s_logisimBus26[3:0]),
.muxIn_1(s_logisimBus56[3:0]),
.muxOut(s_logisimBus16[3:0]),
.sel(s_logisimNet28));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_12
(.enable(1'b1),
.muxIn_0(s_logisimBus16[3:0]),
.muxIn_1(s_logisimBus57[3:0]),
.muxOut(s_logisimBus18[3:0]),
.sel(s_logisimNet20));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_13
(.enable(1'b1),
.muxIn_0(s_logisimBus18[3:0]),
.muxIn_1(s_logisimBus58[3:0]),
.muxOut(s_logisimBus38[3:0]),
.sel(s_logisimNet0));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_14
(.enable(1'b1),
.muxIn_0(s_logisimBus38[3:0]),
.muxIn_1(s_logisimBus59[3:0]),
.muxOut(s_logisimBus24[3:0]),
.sel(s_logisimNet41));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_15
(.enable(1'b1),
.muxIn_0(s_logisimBus24[3:0]),
.muxIn_1(s_logisimBus60[3:0]),
.muxOut(s_logisimBus7[3:0]),
.sel(s_logisimNet19));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_16
(.enable(1'b1),
.muxIn_0(s_logisimBus7[3:0]),
.muxIn_1(s_logisimBus61[3:0]),
.muxOut(s_logisimBus33[3:0]),
.sel(s_logisimNet1));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_17
(.enable(1'b1),
.muxIn_0(s_logisimBus33[3:0]),
.muxIn_1(s_logisimBus62[3:0]),
.muxOut(s_logisimBus8[3:0]),
.sel(s_logisimNet27));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_18
(.enable(1'b1),
.muxIn_0(s_logisimBus8[3:0]),
.muxIn_1(s_logisimBus63[3:0]),
.muxOut(s_logisimBus34[3:0]),
.sel(s_logisimNet42));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_19
(.enable(1'b1),
.muxIn_0(s_logisimBus34[3:0]),
.muxIn_1(s_logisimBus64[3:0]),
.muxOut(s_logisimBus10[3:0]),
.sel(s_logisimNet29));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_20
(.enable(1'b1),
.muxIn_0(s_logisimBus10[3:0]),
.muxIn_1(s_logisimBus65[3:0]),
.muxOut(s_logisimBus35[3:0]),
.sel(s_logisimNet43));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_21
(.enable(1'b1),
.muxIn_0(s_logisimBus35[3:0]),
.muxIn_1(s_logisimBus66[3:0]),
.muxOut(s_logisimBus11[3:0]),
.sel(s_logisimNet36));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_22
(.enable(1'b1),
.muxIn_0(s_logisimBus11[3:0]),
.muxIn_1(s_logisimBus67[3:0]),
.muxOut(s_logisimBus25[3:0]),
.sel(s_logisimNet6));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_23
(.enable(1'b1),
.muxIn_0(s_logisimBus25[3:0]),
.muxIn_1(s_logisimBus68[3:0]),
.muxOut(s_logisimBus39[3:0]),
.sel(s_logisimNet44));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_24
(.enable(1'b1),
.muxIn_0(s_logisimBus39[3:0]),
.muxIn_1(s_logisimBus69[3:0]),
.muxOut(s_logisimBus30[3:0]),
.sel(s_logisimNet45));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_25
(.aEqualsB(s_logisimNet71),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus70[5:0]),
.dataB(s_logisimBus15[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_26
(.aEqualsB(s_logisimNet4),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus72[5:0]),
.dataB(s_logisimBus15[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_27
(.aEqualsB(s_logisimNet5),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus73[5:0]),
.dataB(s_logisimBus15[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_28
(.aEqualsB(s_logisimNet12),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus74[5:0]),
.dataB(s_logisimBus15[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_29
(.aEqualsB(s_logisimNet21),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus75[5:0]),
.dataB(s_logisimBus15[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_30
(.aEqualsB(s_logisimNet2),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus76[5:0]),
.dataB(s_logisimBus15[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_31
(.aEqualsB(s_logisimNet32),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus77[5:0]),
.dataB(s_logisimBus15[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_32
(.aEqualsB(s_logisimNet28),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus78[5:0]),
.dataB(s_logisimBus15[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_33
(.aEqualsB(s_logisimNet20),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus79[5:0]),
.dataB(s_logisimBus15[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_34
(.aEqualsB(s_logisimNet0),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus80[5:0]),
.dataB(s_logisimBus15[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_35
(.aEqualsB(s_logisimNet41),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus81[5:0]),
.dataB(s_logisimBus15[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_36
(.aEqualsB(s_logisimNet19),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus82[5:0]),
.dataB(s_logisimBus15[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_37
(.aEqualsB(s_logisimNet1),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus83[5:0]),
.dataB(s_logisimBus15[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_38
(.aEqualsB(s_logisimNet46),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus84[5:0]),
.dataB(s_logisimBus15[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_39
(.aEqualsB(s_logisimNet31),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus85[5:0]),
.dataB(s_logisimBus9[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_40
(.aEqualsB(s_logisimNet27),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus86[5:0]),
.dataB(s_logisimBus9[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_41
(.aEqualsB(s_logisimNet42),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus87[5:0]),
.dataB(s_logisimBus9[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_42
(.aEqualsB(s_logisimNet29),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus88[5:0]),
.dataB(s_logisimBus9[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_43
(.aEqualsB(s_logisimNet43),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus89[5:0]),
.dataB(s_logisimBus9[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_44
(.aEqualsB(s_logisimNet36),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus90[5:0]),
.dataB(s_logisimBus9[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_45
(.aEqualsB(s_logisimNet6),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus91[5:0]),
.dataB(s_logisimBus9[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_46
(.aEqualsB(s_logisimNet22),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus92[5:0]),
.dataB(s_logisimBus9[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_47
(.aEqualsB(s_logisimNet44),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus93[5:0]),
.dataB(s_logisimBus9[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_48
(.aEqualsB(s_logisimNet3),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus94[5:0]),
.dataB(s_logisimBus9[5:0]));
endmodule