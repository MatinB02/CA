/******************************************************************************
 ** Logisim-evolution goes FPGA automatic generated Verilog code             **
 ** https://github.com/logisim-evolution/                                    **
 **                                                                          **
 ** Component : fadd                                                         **
 **                                                                          **
 *****************************************************************************/

module fadd( INFINITY_PIN,
             NAN_PIN,
             a,
             b,
             res );

   /*******************************************************************************
   ** The inputs are defined here                                                **
   *******************************************************************************/
   input [31:0] a;
   input [31:0] b;

   /*******************************************************************************
   ** The outputs are defined here                                               **
   *******************************************************************************/
   output        INFINITY_PIN;
   output        NAN_PIN;
   output [31:0] res;

   /*******************************************************************************
   ** The wires are defined here                                                 **
   *******************************************************************************/
   wire [31:0] s_logisimBus1;
   wire [22:0] s_logisimBus100;
   wire [22:0] s_logisimBus101;
   wire [31:0] s_logisimBus103;
   wire [22:0] s_logisimBus104;
   wire [31:0] s_logisimBus106;
   wire [8:0]  s_logisimBus107;
   wire [22:0] s_logisimBus108;
   wire [1:0]  s_logisimBus109;
   wire [31:0] s_logisimBus11;
   wire [31:0] s_logisimBus110;
   wire [22:0] s_logisimBus114;
   wire [31:0] s_logisimBus115;
   wire [22:0] s_logisimBus117;
   wire [7:0]  s_logisimBus119;
   wire [22:0] s_logisimBus12;
   wire [22:0] s_logisimBus123;
   wire [22:0] s_logisimBus126;
   wire [31:0] s_logisimBus127;
   wire [22:0] s_logisimBus128;
   wire [1:0]  s_logisimBus13;
   wire [8:0]  s_logisimBus131;
   wire [31:0] s_logisimBus132;
   wire [31:0] s_logisimBus133;
   wire [31:0] s_logisimBus134;
   wire [22:0] s_logisimBus135;
   wire [7:0]  s_logisimBus136;
   wire [7:0]  s_logisimBus137;
   wire [8:0]  s_logisimBus14;
   wire [7:0]  s_logisimBus140;
   wire [21:0] s_logisimBus141;
   wire [22:0] s_logisimBus142;
   wire [31:0] s_logisimBus144;
   wire [31:0] s_logisimBus146;
   wire [22:0] s_logisimBus147;
   wire [22:0] s_logisimBus148;
   wire [22:0] s_logisimBus149;
   wire [7:0]  s_logisimBus150;
   wire [7:0]  s_logisimBus151;
   wire [31:0] s_logisimBus153;
   wire [22:0] s_logisimBus20;
   wire [8:0]  s_logisimBus22;
   wire [31:0] s_logisimBus23;
   wire [31:0] s_logisimBus24;
   wire [23:0] s_logisimBus27;
   wire [8:0]  s_logisimBus29;
   wire [22:0] s_logisimBus3;
   wire [31:0] s_logisimBus32;
   wire [4:0]  s_logisimBus33;
   wire [22:0] s_logisimBus34;
   wire [8:0]  s_logisimBus35;
   wire [7:0]  s_logisimBus36;
   wire [7:0]  s_logisimBus37;
   wire [23:0] s_logisimBus4;
   wire [31:0] s_logisimBus42;
   wire [1:0]  s_logisimBus43;
   wire [63:0] s_logisimBus47;
   wire [8:0]  s_logisimBus48;
   wire [7:0]  s_logisimBus49;
   wire [8:0]  s_logisimBus5;
   wire [22:0] s_logisimBus50;
   wire [31:0] s_logisimBus52;
   wire [31:0] s_logisimBus53;
   wire [31:0] s_logisimBus57;
   wire [22:0] s_logisimBus58;
   wire [7:0]  s_logisimBus6;
   wire [8:0]  s_logisimBus60;
   wire [31:0] s_logisimBus61;
   wire [22:0] s_logisimBus68;
   wire [8:0]  s_logisimBus69;
   wire [31:0] s_logisimBus75;
   wire [31:0] s_logisimBus78;
   wire [31:0] s_logisimBus80;
   wire [63:0] s_logisimBus82;
   wire [22:0] s_logisimBus83;
   wire [7:0]  s_logisimBus84;
   wire [22:0] s_logisimBus85;
   wire [8:0]  s_logisimBus87;
   wire [8:0]  s_logisimBus88;
   wire [31:0] s_logisimBus89;
   wire [31:0] s_logisimBus9;
   wire [4:0]  s_logisimBus91;
   wire [7:0]  s_logisimBus93;
   wire [31:0] s_logisimBus94;
   wire [7:0]  s_logisimBus97;
   wire        s_logisimNet0;
   wire        s_logisimNet10;
   wire        s_logisimNet102;
   wire        s_logisimNet105;
   wire        s_logisimNet111;
   wire        s_logisimNet112;
   wire        s_logisimNet116;
   wire        s_logisimNet118;
   wire        s_logisimNet120;
   wire        s_logisimNet121;
   wire        s_logisimNet122;
   wire        s_logisimNet124;
   wire        s_logisimNet125;
   wire        s_logisimNet129;
   wire        s_logisimNet130;
   wire        s_logisimNet138;
   wire        s_logisimNet139;
   wire        s_logisimNet143;
   wire        s_logisimNet145;
   wire        s_logisimNet15;
   wire        s_logisimNet152;
   wire        s_logisimNet156;
   wire        s_logisimNet157;
   wire        s_logisimNet158;
   wire        s_logisimNet159;
   wire        s_logisimNet16;
   wire        s_logisimNet17;
   wire        s_logisimNet18;
   wire        s_logisimNet19;
   wire        s_logisimNet2;
   wire        s_logisimNet21;
   wire        s_logisimNet25;
   wire        s_logisimNet26;
   wire        s_logisimNet28;
   wire        s_logisimNet30;
   wire        s_logisimNet38;
   wire        s_logisimNet40;
   wire        s_logisimNet41;
   wire        s_logisimNet44;
   wire        s_logisimNet45;
   wire        s_logisimNet46;
   wire        s_logisimNet51;
   wire        s_logisimNet55;
   wire        s_logisimNet56;
   wire        s_logisimNet59;
   wire        s_logisimNet62;
   wire        s_logisimNet63;
   wire        s_logisimNet64;
   wire        s_logisimNet65;
   wire        s_logisimNet66;
   wire        s_logisimNet67;
   wire        s_logisimNet7;
   wire        s_logisimNet70;
   wire        s_logisimNet71;
   wire        s_logisimNet72;
   wire        s_logisimNet73;
   wire        s_logisimNet74;
   wire        s_logisimNet76;
   wire        s_logisimNet77;
   wire        s_logisimNet79;
   wire        s_logisimNet8;
   wire        s_logisimNet81;
   wire        s_logisimNet90;
   wire        s_logisimNet92;
   wire        s_logisimNet95;
   wire        s_logisimNet96;
   wire        s_logisimNet99;

   /*******************************************************************************
   ** The module functionality is described here                                 **
   *******************************************************************************/

   /*******************************************************************************
   ** Here all wiring is defined                                                 **
   *******************************************************************************/
   assign s_logisimBus101[0]  = s_logisimBus141[0];
   assign s_logisimBus101[10] = s_logisimBus141[10];
   assign s_logisimBus101[11] = s_logisimBus141[11];
   assign s_logisimBus101[12] = s_logisimBus141[12];
   assign s_logisimBus101[13] = s_logisimBus141[13];
   assign s_logisimBus101[14] = s_logisimBus141[14];
   assign s_logisimBus101[15] = s_logisimBus141[15];
   assign s_logisimBus101[16] = s_logisimBus141[16];
   assign s_logisimBus101[17] = s_logisimBus141[17];
   assign s_logisimBus101[18] = s_logisimBus141[18];
   assign s_logisimBus101[19] = s_logisimBus141[19];
   assign s_logisimBus101[1]  = s_logisimBus141[1];
   assign s_logisimBus101[20] = s_logisimBus141[20];
   assign s_logisimBus101[21] = s_logisimBus141[21];
   assign s_logisimBus101[22] = s_logisimNet72;
   assign s_logisimBus101[2]  = s_logisimBus141[2];
   assign s_logisimBus101[3]  = s_logisimBus141[3];
   assign s_logisimBus101[4]  = s_logisimBus141[4];
   assign s_logisimBus101[5]  = s_logisimBus141[5];
   assign s_logisimBus101[6]  = s_logisimBus141[6];
   assign s_logisimBus101[7]  = s_logisimBus141[7];
   assign s_logisimBus101[8]  = s_logisimBus141[8];
   assign s_logisimBus101[9]  = s_logisimBus141[9];
   assign s_logisimBus135[0]  = s_logisimBus127[0];
   assign s_logisimBus135[10] = s_logisimBus127[10];
   assign s_logisimBus135[11] = s_logisimBus127[11];
   assign s_logisimBus135[12] = s_logisimBus127[12];
   assign s_logisimBus135[13] = s_logisimBus127[13];
   assign s_logisimBus135[14] = s_logisimBus127[14];
   assign s_logisimBus135[15] = s_logisimBus127[15];
   assign s_logisimBus135[16] = s_logisimBus127[16];
   assign s_logisimBus135[17] = s_logisimBus127[17];
   assign s_logisimBus135[18] = s_logisimBus127[18];
   assign s_logisimBus135[19] = s_logisimBus127[19];
   assign s_logisimBus135[1]  = s_logisimBus127[1];
   assign s_logisimBus135[20] = s_logisimBus127[20];
   assign s_logisimBus135[21] = s_logisimBus127[21];
   assign s_logisimBus135[22] = s_logisimBus127[22];
   assign s_logisimBus135[2]  = s_logisimBus127[2];
   assign s_logisimBus135[3]  = s_logisimBus127[3];
   assign s_logisimBus135[4]  = s_logisimBus127[4];
   assign s_logisimBus135[5]  = s_logisimBus127[5];
   assign s_logisimBus135[6]  = s_logisimBus127[6];
   assign s_logisimBus135[7]  = s_logisimBus127[7];
   assign s_logisimBus135[8]  = s_logisimBus127[8];
   assign s_logisimBus135[9]  = s_logisimBus127[9];
   assign s_logisimBus140[0]  = s_logisimBus134[23];
   assign s_logisimBus140[1]  = s_logisimBus134[24];
   assign s_logisimBus140[2]  = s_logisimBus134[25];
   assign s_logisimBus140[3]  = s_logisimBus134[26];
   assign s_logisimBus140[4]  = s_logisimBus134[27];
   assign s_logisimBus140[5]  = s_logisimBus134[28];
   assign s_logisimBus140[6]  = s_logisimBus134[29];
   assign s_logisimBus140[7]  = s_logisimBus134[30];
   assign s_logisimBus141[0]  = s_logisimBus149[1];
   assign s_logisimBus141[10] = s_logisimBus149[11];
   assign s_logisimBus141[11] = s_logisimBus149[12];
   assign s_logisimBus141[12] = s_logisimBus149[13];
   assign s_logisimBus141[13] = s_logisimBus149[14];
   assign s_logisimBus141[14] = s_logisimBus149[15];
   assign s_logisimBus141[15] = s_logisimBus149[16];
   assign s_logisimBus141[16] = s_logisimBus149[17];
   assign s_logisimBus141[17] = s_logisimBus149[18];
   assign s_logisimBus141[18] = s_logisimBus149[19];
   assign s_logisimBus141[19] = s_logisimBus149[20];
   assign s_logisimBus141[1]  = s_logisimBus149[2];
   assign s_logisimBus141[20] = s_logisimBus149[21];
   assign s_logisimBus141[21] = s_logisimBus149[22];
   assign s_logisimBus141[2]  = s_logisimBus149[3];
   assign s_logisimBus141[3]  = s_logisimBus149[4];
   assign s_logisimBus141[4]  = s_logisimBus149[5];
   assign s_logisimBus141[5]  = s_logisimBus149[6];
   assign s_logisimBus141[6]  = s_logisimBus149[7];
   assign s_logisimBus141[7]  = s_logisimBus149[8];
   assign s_logisimBus141[8]  = s_logisimBus149[9];
   assign s_logisimBus141[9]  = s_logisimBus149[10];
   assign s_logisimBus148[0]  = s_logisimBus134[0];
   assign s_logisimBus148[10] = s_logisimBus134[10];
   assign s_logisimBus148[11] = s_logisimBus134[11];
   assign s_logisimBus148[12] = s_logisimBus134[12];
   assign s_logisimBus148[13] = s_logisimBus134[13];
   assign s_logisimBus148[14] = s_logisimBus134[14];
   assign s_logisimBus148[15] = s_logisimBus134[15];
   assign s_logisimBus148[16] = s_logisimBus134[16];
   assign s_logisimBus148[17] = s_logisimBus134[17];
   assign s_logisimBus148[18] = s_logisimBus134[18];
   assign s_logisimBus148[19] = s_logisimBus134[19];
   assign s_logisimBus148[1]  = s_logisimBus134[1];
   assign s_logisimBus148[20] = s_logisimBus134[20];
   assign s_logisimBus148[21] = s_logisimBus134[21];
   assign s_logisimBus148[22] = s_logisimBus134[22];
   assign s_logisimBus148[2]  = s_logisimBus134[2];
   assign s_logisimBus148[3]  = s_logisimBus134[3];
   assign s_logisimBus148[4]  = s_logisimBus134[4];
   assign s_logisimBus148[5]  = s_logisimBus134[5];
   assign s_logisimBus148[6]  = s_logisimBus134[6];
   assign s_logisimBus148[7]  = s_logisimBus134[7];
   assign s_logisimBus148[8]  = s_logisimBus134[8];
   assign s_logisimBus148[9]  = s_logisimBus134[9];
   assign s_logisimBus151[0]  = s_logisimBus127[23];
   assign s_logisimBus151[1]  = s_logisimBus127[24];
   assign s_logisimBus151[2]  = s_logisimBus127[25];
   assign s_logisimBus151[3]  = s_logisimBus127[26];
   assign s_logisimBus151[4]  = s_logisimBus127[27];
   assign s_logisimBus151[5]  = s_logisimBus127[28];
   assign s_logisimBus151[6]  = s_logisimBus127[29];
   assign s_logisimBus151[7]  = s_logisimBus127[30];
   assign s_logisimBus22[0]   = s_logisimBus140[0];
   assign s_logisimBus22[1]   = s_logisimBus140[1];
   assign s_logisimBus22[2]   = s_logisimBus140[2];
   assign s_logisimBus22[3]   = s_logisimBus140[3];
   assign s_logisimBus22[4]   = s_logisimBus140[4];
   assign s_logisimBus22[5]   = s_logisimBus140[5];
   assign s_logisimBus22[6]   = s_logisimBus140[6];
   assign s_logisimBus22[7]   = s_logisimBus140[7];
   assign s_logisimBus27[0]   = s_logisimBus148[0];
   assign s_logisimBus27[10]  = s_logisimBus148[10];
   assign s_logisimBus27[11]  = s_logisimBus148[11];
   assign s_logisimBus27[12]  = s_logisimBus148[12];
   assign s_logisimBus27[13]  = s_logisimBus148[13];
   assign s_logisimBus27[14]  = s_logisimBus148[14];
   assign s_logisimBus27[15]  = s_logisimBus148[15];
   assign s_logisimBus27[16]  = s_logisimBus148[16];
   assign s_logisimBus27[17]  = s_logisimBus148[17];
   assign s_logisimBus27[18]  = s_logisimBus148[18];
   assign s_logisimBus27[19]  = s_logisimBus148[19];
   assign s_logisimBus27[1]   = s_logisimBus148[1];
   assign s_logisimBus27[20]  = s_logisimBus148[20];
   assign s_logisimBus27[21]  = s_logisimBus148[21];
   assign s_logisimBus27[22]  = s_logisimBus148[22];
   assign s_logisimBus27[2]   = s_logisimBus148[2];
   assign s_logisimBus27[3]   = s_logisimBus148[3];
   assign s_logisimBus27[4]   = s_logisimBus148[4];
   assign s_logisimBus27[5]   = s_logisimBus148[5];
   assign s_logisimBus27[6]   = s_logisimBus148[6];
   assign s_logisimBus27[7]   = s_logisimBus148[7];
   assign s_logisimBus27[8]   = s_logisimBus148[8];
   assign s_logisimBus27[9]   = s_logisimBus148[9];
   assign s_logisimBus29[0]   = s_logisimBus140[0];
   assign s_logisimBus29[1]   = s_logisimBus140[1];
   assign s_logisimBus29[2]   = s_logisimBus140[2];
   assign s_logisimBus29[3]   = s_logisimBus140[3];
   assign s_logisimBus29[4]   = s_logisimBus140[4];
   assign s_logisimBus29[5]   = s_logisimBus140[5];
   assign s_logisimBus29[6]   = s_logisimBus140[6];
   assign s_logisimBus29[7]   = s_logisimBus140[7];
   assign s_logisimBus32[31]  = s_logisimNet156;
   assign s_logisimBus35[0]   = s_logisimBus151[0];
   assign s_logisimBus35[1]   = s_logisimBus151[1];
   assign s_logisimBus35[2]   = s_logisimBus151[2];
   assign s_logisimBus35[3]   = s_logisimBus151[3];
   assign s_logisimBus35[4]   = s_logisimBus151[4];
   assign s_logisimBus35[5]   = s_logisimBus151[5];
   assign s_logisimBus35[6]   = s_logisimBus151[6];
   assign s_logisimBus35[7]   = s_logisimBus151[7];
   assign s_logisimBus48[0]   = s_logisimBus140[0];
   assign s_logisimBus48[1]   = s_logisimBus140[1];
   assign s_logisimBus48[2]   = s_logisimBus140[2];
   assign s_logisimBus48[3]   = s_logisimBus140[3];
   assign s_logisimBus48[4]   = s_logisimBus140[4];
   assign s_logisimBus48[5]   = s_logisimBus140[5];
   assign s_logisimBus48[6]   = s_logisimBus140[6];
   assign s_logisimBus48[7]   = s_logisimBus140[7];
   assign s_logisimBus4[0]    = s_logisimBus135[0];
   assign s_logisimBus4[10]   = s_logisimBus135[10];
   assign s_logisimBus4[11]   = s_logisimBus135[11];
   assign s_logisimBus4[12]   = s_logisimBus135[12];
   assign s_logisimBus4[13]   = s_logisimBus135[13];
   assign s_logisimBus4[14]   = s_logisimBus135[14];
   assign s_logisimBus4[15]   = s_logisimBus135[15];
   assign s_logisimBus4[16]   = s_logisimBus135[16];
   assign s_logisimBus4[17]   = s_logisimBus135[17];
   assign s_logisimBus4[18]   = s_logisimBus135[18];
   assign s_logisimBus4[19]   = s_logisimBus135[19];
   assign s_logisimBus4[1]    = s_logisimBus135[1];
   assign s_logisimBus4[20]   = s_logisimBus135[20];
   assign s_logisimBus4[21]   = s_logisimBus135[21];
   assign s_logisimBus4[22]   = s_logisimBus135[22];
   assign s_logisimBus4[2]    = s_logisimBus135[2];
   assign s_logisimBus4[3]    = s_logisimBus135[3];
   assign s_logisimBus4[4]    = s_logisimBus135[4];
   assign s_logisimBus4[5]    = s_logisimBus135[5];
   assign s_logisimBus4[6]    = s_logisimBus135[6];
   assign s_logisimBus4[7]    = s_logisimBus135[7];
   assign s_logisimBus4[8]    = s_logisimBus135[8];
   assign s_logisimBus4[9]    = s_logisimBus135[9];
   assign s_logisimBus5[0]    = s_logisimBus151[0];
   assign s_logisimBus5[1]    = s_logisimBus151[1];
   assign s_logisimBus5[2]    = s_logisimBus151[2];
   assign s_logisimBus5[3]    = s_logisimBus151[3];
   assign s_logisimBus5[4]    = s_logisimBus151[4];
   assign s_logisimBus5[5]    = s_logisimBus151[5];
   assign s_logisimBus5[6]    = s_logisimBus151[6];
   assign s_logisimBus5[7]    = s_logisimBus151[7];
   assign s_logisimBus69[0]   = s_logisimBus151[0];
   assign s_logisimBus69[1]   = s_logisimBus151[1];
   assign s_logisimBus69[2]   = s_logisimBus151[2];
   assign s_logisimBus69[3]   = s_logisimBus151[3];
   assign s_logisimBus69[4]   = s_logisimBus151[4];
   assign s_logisimBus69[5]   = s_logisimBus151[5];
   assign s_logisimBus69[6]   = s_logisimBus151[6];
   assign s_logisimBus69[7]   = s_logisimBus151[7];
   assign s_logisimBus87[0]   = s_logisimBus140[0];
   assign s_logisimBus87[1]   = s_logisimBus140[1];
   assign s_logisimBus87[2]   = s_logisimBus140[2];
   assign s_logisimBus87[3]   = s_logisimBus140[3];
   assign s_logisimBus87[4]   = s_logisimBus140[4];
   assign s_logisimBus87[5]   = s_logisimBus140[5];
   assign s_logisimBus87[6]   = s_logisimBus140[6];
   assign s_logisimBus87[7]   = s_logisimBus140[7];
   assign s_logisimBus88[0]   = s_logisimBus151[0];
   assign s_logisimBus88[1]   = s_logisimBus151[1];
   assign s_logisimBus88[2]   = s_logisimBus151[2];
   assign s_logisimBus88[3]   = s_logisimBus151[3];
   assign s_logisimBus88[4]   = s_logisimBus151[4];
   assign s_logisimBus88[5]   = s_logisimBus151[5];
   assign s_logisimBus88[6]   = s_logisimBus151[6];
   assign s_logisimBus88[7]   = s_logisimBus151[7];
   assign s_logisimNet156     = s_logisimBus127[31];
   assign s_logisimNet72      = s_logisimBus43[0];

   /*******************************************************************************
   ** Here all input connections are defined                                     **
   *******************************************************************************/
   assign s_logisimBus127[31:0] = a;
   assign s_logisimBus134[31:0] = b;

   /*******************************************************************************
   ** Here all output connections are defined                                    **
   *******************************************************************************/
   assign INFINITY_PIN = s_logisimNet105;
   assign NAN_PIN      = s_logisimNet129;
   assign res          = s_logisimBus24[31:0];

   /*******************************************************************************
   ** Here all in-lined components are defined                                   **
   *******************************************************************************/

   // Constant
   assign  s_logisimBus146[31:0]  =  32'h00000019;


   // Constant
   assign  s_logisimBus35[8]  =  1'b0;


   // Constant
   assign  s_logisimBus48[8]  =  1'b0;


   // Constant
   assign  s_logisimBus91[4:0]  =  {1'b0, 4'h1};


   // Constant
   assign  s_logisimBus22[8]  =  1'b0;


   // Constant
   assign  s_logisimBus69[8]  =  1'b0;


   // Constant
   assign  s_logisimBus33[4:0]  =  {1'b0, 4'h1};


   // Constant
   assign  s_logisimNet118  =  1'b0;


   // Constant
   assign  s_logisimBus75[31:0]  =  32'h00000019;


   // Constant
   assign  s_logisimNet46  =  1'b0;


   // Constant
   assign  s_logisimBus131[8:0]  =  {1'b0, 8'hC0};


   // Constant
   assign  s_logisimBus107[8:0]  =  {1'b0, 8'hC0};


   // Constant
   assign  s_logisimBus110[31:0]  =  32'h00000001;


   // Constant
   assign  s_logisimBus128[22:0]  =  {3'b000, 20'h00001};


   // Constant
   assign  s_logisimBus153[31:0]  =  32'h00000001;


   // Constant
   assign  s_logisimBus104[22:0]  =  {3'b000, 20'h00001};


   // Constant
   assign  s_logisimBus37[7:0]  =  8'hFF;


   // Constant
   assign  s_logisimBus114[22:0]  =  {3'b000, 20'h00000};


   // Constant
   assign  s_logisimBus136[7:0]  =  8'hFF;


   // Constant
   assign  s_logisimBus85[22:0]  =  {3'b000, 20'h00000};


   // Constant
   assign  s_logisimBus109[1:0]  =  2'b10;


   // Constant
   assign  s_logisimBus84[7:0]  =  8'hFF;


   // Constant
   assign  s_logisimBus12[22:0]  =  {3'b000, 20'h00000};


   // Constant
   assign  s_logisimBus49[7:0]  =  8'hFF;


   // Constant
   assign  s_logisimBus123[22:0]  =  {3'b000, 20'h00000};


   // Bit Extender
   assign  s_logisimBus1[0]  =  s_logisimBus97[0];
   assign  s_logisimBus1[1]  =  s_logisimBus97[1];
   assign  s_logisimBus1[2]  =  s_logisimBus97[2];
   assign  s_logisimBus1[3]  =  s_logisimBus97[3];
   assign  s_logisimBus1[4]  =  s_logisimBus97[4];
   assign  s_logisimBus1[5]  =  s_logisimBus97[5];
   assign  s_logisimBus1[6]  =  s_logisimBus97[6];
   assign  s_logisimBus1[7]  =  s_logisimBus97[7];
   assign  s_logisimBus1[8]  =  1'b0;
   assign  s_logisimBus1[9]  =  1'b0;
   assign  s_logisimBus1[10]  =  1'b0;
   assign  s_logisimBus1[11]  =  1'b0;
   assign  s_logisimBus1[12]  =  1'b0;
   assign  s_logisimBus1[13]  =  1'b0;
   assign  s_logisimBus1[14]  =  1'b0;
   assign  s_logisimBus1[15]  =  1'b0;
   assign  s_logisimBus1[16]  =  1'b0;
   assign  s_logisimBus1[17]  =  1'b0;
   assign  s_logisimBus1[18]  =  1'b0;
   assign  s_logisimBus1[19]  =  1'b0;
   assign  s_logisimBus1[20]  =  1'b0;
   assign  s_logisimBus1[21]  =  1'b0;
   assign  s_logisimBus1[22]  =  1'b0;
   assign  s_logisimBus1[23]  =  1'b0;
   assign  s_logisimBus1[24]  =  1'b0;
   assign  s_logisimBus1[25]  =  1'b0;
   assign  s_logisimBus1[26]  =  1'b0;
   assign  s_logisimBus1[27]  =  1'b0;
   assign  s_logisimBus1[28]  =  1'b0;
   assign  s_logisimBus1[29]  =  1'b0;
   assign  s_logisimBus1[30]  =  1'b0;
   assign  s_logisimBus1[31]  =  1'b0;


   // Bit Extender
   assign  s_logisimBus53[0]  =  s_logisimBus137[0];
   assign  s_logisimBus53[1]  =  s_logisimBus137[1];
   assign  s_logisimBus53[2]  =  s_logisimBus137[2];
   assign  s_logisimBus53[3]  =  s_logisimBus137[3];
   assign  s_logisimBus53[4]  =  s_logisimBus137[4];
   assign  s_logisimBus53[5]  =  s_logisimBus137[5];
   assign  s_logisimBus53[6]  =  s_logisimBus137[6];
   assign  s_logisimBus53[7]  =  s_logisimBus137[7];
   assign  s_logisimBus53[8]  =  1'b0;
   assign  s_logisimBus53[9]  =  1'b0;
   assign  s_logisimBus53[10]  =  1'b0;
   assign  s_logisimBus53[11]  =  1'b0;
   assign  s_logisimBus53[12]  =  1'b0;
   assign  s_logisimBus53[13]  =  1'b0;
   assign  s_logisimBus53[14]  =  1'b0;
   assign  s_logisimBus53[15]  =  1'b0;
   assign  s_logisimBus53[16]  =  1'b0;
   assign  s_logisimBus53[17]  =  1'b0;
   assign  s_logisimBus53[18]  =  1'b0;
   assign  s_logisimBus53[19]  =  1'b0;
   assign  s_logisimBus53[20]  =  1'b0;
   assign  s_logisimBus53[21]  =  1'b0;
   assign  s_logisimBus53[22]  =  1'b0;
   assign  s_logisimBus53[23]  =  1'b0;
   assign  s_logisimBus53[24]  =  1'b0;
   assign  s_logisimBus53[25]  =  1'b0;
   assign  s_logisimBus53[26]  =  1'b0;
   assign  s_logisimBus53[27]  =  1'b0;
   assign  s_logisimBus53[28]  =  1'b0;
   assign  s_logisimBus53[29]  =  1'b0;
   assign  s_logisimBus53[30]  =  1'b0;
   assign  s_logisimBus53[31]  =  1'b0;


   // Constant
   assign  s_logisimBus150[7:0]  =  8'h00;


   // Bit Extender
   assign  s_logisimBus13[0]  =  s_logisimNet124;
   assign  s_logisimBus13[1]  =  1'b0;


   // Constant
   assign  s_logisimBus93[7:0]  =  8'h00;


   // Bit Extender
   assign  s_logisimBus9[0]  =  s_logisimBus4[0];
   assign  s_logisimBus9[1]  =  s_logisimBus4[1];
   assign  s_logisimBus9[2]  =  s_logisimBus4[2];
   assign  s_logisimBus9[3]  =  s_logisimBus4[3];
   assign  s_logisimBus9[4]  =  s_logisimBus4[4];
   assign  s_logisimBus9[5]  =  s_logisimBus4[5];
   assign  s_logisimBus9[6]  =  s_logisimBus4[6];
   assign  s_logisimBus9[7]  =  s_logisimBus4[7];
   assign  s_logisimBus9[8]  =  s_logisimBus4[8];
   assign  s_logisimBus9[9]  =  s_logisimBus4[9];
   assign  s_logisimBus9[10]  =  s_logisimBus4[10];
   assign  s_logisimBus9[11]  =  s_logisimBus4[11];
   assign  s_logisimBus9[12]  =  s_logisimBus4[12];
   assign  s_logisimBus9[13]  =  s_logisimBus4[13];
   assign  s_logisimBus9[14]  =  s_logisimBus4[14];
   assign  s_logisimBus9[15]  =  s_logisimBus4[15];
   assign  s_logisimBus9[16]  =  s_logisimBus4[16];
   assign  s_logisimBus9[17]  =  s_logisimBus4[17];
   assign  s_logisimBus9[18]  =  s_logisimBus4[18];
   assign  s_logisimBus9[19]  =  s_logisimBus4[19];
   assign  s_logisimBus9[20]  =  s_logisimBus4[20];
   assign  s_logisimBus9[21]  =  s_logisimBus4[21];
   assign  s_logisimBus9[22]  =  s_logisimBus4[22];
   assign  s_logisimBus9[23]  =  s_logisimBus4[23];
   assign  s_logisimBus9[24]  =  1'b0;
   assign  s_logisimBus9[25]  =  1'b0;
   assign  s_logisimBus9[26]  =  1'b0;
   assign  s_logisimBus9[27]  =  1'b0;
   assign  s_logisimBus9[28]  =  1'b0;
   assign  s_logisimBus9[29]  =  1'b0;
   assign  s_logisimBus9[30]  =  1'b0;
   assign  s_logisimBus9[31]  =  1'b0;


   // Bit Extender
   assign  s_logisimBus11[0]  =  s_logisimBus27[0];
   assign  s_logisimBus11[1]  =  s_logisimBus27[1];
   assign  s_logisimBus11[2]  =  s_logisimBus27[2];
   assign  s_logisimBus11[3]  =  s_logisimBus27[3];
   assign  s_logisimBus11[4]  =  s_logisimBus27[4];
   assign  s_logisimBus11[5]  =  s_logisimBus27[5];
   assign  s_logisimBus11[6]  =  s_logisimBus27[6];
   assign  s_logisimBus11[7]  =  s_logisimBus27[7];
   assign  s_logisimBus11[8]  =  s_logisimBus27[8];
   assign  s_logisimBus11[9]  =  s_logisimBus27[9];
   assign  s_logisimBus11[10]  =  s_logisimBus27[10];
   assign  s_logisimBus11[11]  =  s_logisimBus27[11];
   assign  s_logisimBus11[12]  =  s_logisimBus27[12];
   assign  s_logisimBus11[13]  =  s_logisimBus27[13];
   assign  s_logisimBus11[14]  =  s_logisimBus27[14];
   assign  s_logisimBus11[15]  =  s_logisimBus27[15];
   assign  s_logisimBus11[16]  =  s_logisimBus27[16];
   assign  s_logisimBus11[17]  =  s_logisimBus27[17];
   assign  s_logisimBus11[18]  =  s_logisimBus27[18];
   assign  s_logisimBus11[19]  =  s_logisimBus27[19];
   assign  s_logisimBus11[20]  =  s_logisimBus27[20];
   assign  s_logisimBus11[21]  =  s_logisimBus27[21];
   assign  s_logisimBus11[22]  =  s_logisimBus27[22];
   assign  s_logisimBus11[23]  =  s_logisimBus27[23];
   assign  s_logisimBus11[24]  =  1'b0;
   assign  s_logisimBus11[25]  =  1'b0;
   assign  s_logisimBus11[26]  =  1'b0;
   assign  s_logisimBus11[27]  =  1'b0;
   assign  s_logisimBus11[28]  =  1'b0;
   assign  s_logisimBus11[29]  =  1'b0;
   assign  s_logisimBus11[30]  =  1'b0;
   assign  s_logisimBus11[31]  =  1'b0;


   // Constant
   assign  s_logisimNet116  =  1'b1;


   // Constant
   assign  s_logisimNet67  =  1'b0;


   // Constant
   assign  s_logisimNet59  =  1'b1;


   // Constant
   assign  s_logisimNet139  =  1'b0;


   // Constant
   assign  s_logisimBus5[8]  =  1'b0;


   // Constant
   assign  s_logisimBus87[8]  =  1'b0;


   // Constant
   assign  s_logisimBus88[8]  =  1'b0;


   // Constant
   assign  s_logisimBus29[8]  =  1'b0;


   // Bit Extender
   assign  s_logisimBus82[0]  =  s_logisimBus52[0];
   assign  s_logisimBus82[1]  =  s_logisimBus52[1];
   assign  s_logisimBus82[2]  =  s_logisimBus52[2];
   assign  s_logisimBus82[3]  =  s_logisimBus52[3];
   assign  s_logisimBus82[4]  =  s_logisimBus52[4];
   assign  s_logisimBus82[5]  =  s_logisimBus52[5];
   assign  s_logisimBus82[6]  =  s_logisimBus52[6];
   assign  s_logisimBus82[7]  =  s_logisimBus52[7];
   assign  s_logisimBus82[8]  =  s_logisimBus52[8];
   assign  s_logisimBus82[9]  =  s_logisimBus52[9];
   assign  s_logisimBus82[10]  =  s_logisimBus52[10];
   assign  s_logisimBus82[11]  =  s_logisimBus52[11];
   assign  s_logisimBus82[12]  =  s_logisimBus52[12];
   assign  s_logisimBus82[13]  =  s_logisimBus52[13];
   assign  s_logisimBus82[14]  =  s_logisimBus52[14];
   assign  s_logisimBus82[15]  =  s_logisimBus52[15];
   assign  s_logisimBus82[16]  =  s_logisimBus52[16];
   assign  s_logisimBus82[17]  =  s_logisimBus52[17];
   assign  s_logisimBus82[18]  =  s_logisimBus52[18];
   assign  s_logisimBus82[19]  =  s_logisimBus52[19];
   assign  s_logisimBus82[20]  =  s_logisimBus52[20];
   assign  s_logisimBus82[21]  =  s_logisimBus52[21];
   assign  s_logisimBus82[22]  =  s_logisimBus52[22];
   assign  s_logisimBus82[23]  =  s_logisimBus52[23];
   assign  s_logisimBus82[24]  =  s_logisimBus52[24];
   assign  s_logisimBus82[25]  =  s_logisimBus52[25];
   assign  s_logisimBus82[26]  =  s_logisimBus52[26];
   assign  s_logisimBus82[27]  =  s_logisimBus52[27];
   assign  s_logisimBus82[28]  =  s_logisimBus52[28];
   assign  s_logisimBus82[29]  =  s_logisimBus52[29];
   assign  s_logisimBus82[30]  =  s_logisimBus52[30];
   assign  s_logisimBus82[31]  =  s_logisimBus52[31];
   assign  s_logisimBus82[32]  =  1'b0;
   assign  s_logisimBus82[33]  =  1'b0;
   assign  s_logisimBus82[34]  =  1'b0;
   assign  s_logisimBus82[35]  =  1'b0;
   assign  s_logisimBus82[36]  =  1'b0;
   assign  s_logisimBus82[37]  =  1'b0;
   assign  s_logisimBus82[38]  =  1'b0;
   assign  s_logisimBus82[39]  =  1'b0;
   assign  s_logisimBus82[40]  =  1'b0;
   assign  s_logisimBus82[41]  =  1'b0;
   assign  s_logisimBus82[42]  =  1'b0;
   assign  s_logisimBus82[43]  =  1'b0;
   assign  s_logisimBus82[44]  =  1'b0;
   assign  s_logisimBus82[45]  =  1'b0;
   assign  s_logisimBus82[46]  =  1'b0;
   assign  s_logisimBus82[47]  =  1'b0;
   assign  s_logisimBus82[48]  =  1'b0;
   assign  s_logisimBus82[49]  =  1'b0;
   assign  s_logisimBus82[50]  =  1'b0;
   assign  s_logisimBus82[51]  =  1'b0;
   assign  s_logisimBus82[52]  =  1'b0;
   assign  s_logisimBus82[53]  =  1'b0;
   assign  s_logisimBus82[54]  =  1'b0;
   assign  s_logisimBus82[55]  =  1'b0;
   assign  s_logisimBus82[56]  =  1'b0;
   assign  s_logisimBus82[57]  =  1'b0;
   assign  s_logisimBus82[58]  =  1'b0;
   assign  s_logisimBus82[59]  =  1'b0;
   assign  s_logisimBus82[60]  =  1'b0;
   assign  s_logisimBus82[61]  =  1'b0;
   assign  s_logisimBus82[62]  =  1'b0;
   assign  s_logisimBus82[63]  =  1'b0;


   // Bit Extender
   assign  s_logisimBus47[0]  =  s_logisimBus57[0];
   assign  s_logisimBus47[1]  =  s_logisimBus57[1];
   assign  s_logisimBus47[2]  =  s_logisimBus57[2];
   assign  s_logisimBus47[3]  =  s_logisimBus57[3];
   assign  s_logisimBus47[4]  =  s_logisimBus57[4];
   assign  s_logisimBus47[5]  =  s_logisimBus57[5];
   assign  s_logisimBus47[6]  =  s_logisimBus57[6];
   assign  s_logisimBus47[7]  =  s_logisimBus57[7];
   assign  s_logisimBus47[8]  =  s_logisimBus57[8];
   assign  s_logisimBus47[9]  =  s_logisimBus57[9];
   assign  s_logisimBus47[10]  =  s_logisimBus57[10];
   assign  s_logisimBus47[11]  =  s_logisimBus57[11];
   assign  s_logisimBus47[12]  =  s_logisimBus57[12];
   assign  s_logisimBus47[13]  =  s_logisimBus57[13];
   assign  s_logisimBus47[14]  =  s_logisimBus57[14];
   assign  s_logisimBus47[15]  =  s_logisimBus57[15];
   assign  s_logisimBus47[16]  =  s_logisimBus57[16];
   assign  s_logisimBus47[17]  =  s_logisimBus57[17];
   assign  s_logisimBus47[18]  =  s_logisimBus57[18];
   assign  s_logisimBus47[19]  =  s_logisimBus57[19];
   assign  s_logisimBus47[20]  =  s_logisimBus57[20];
   assign  s_logisimBus47[21]  =  s_logisimBus57[21];
   assign  s_logisimBus47[22]  =  s_logisimBus57[22];
   assign  s_logisimBus47[23]  =  s_logisimBus57[23];
   assign  s_logisimBus47[24]  =  s_logisimBus57[24];
   assign  s_logisimBus47[25]  =  s_logisimBus57[25];
   assign  s_logisimBus47[26]  =  s_logisimBus57[26];
   assign  s_logisimBus47[27]  =  s_logisimBus57[27];
   assign  s_logisimBus47[28]  =  s_logisimBus57[28];
   assign  s_logisimBus47[29]  =  s_logisimBus57[29];
   assign  s_logisimBus47[30]  =  s_logisimBus57[30];
   assign  s_logisimBus47[31]  =  s_logisimBus57[31];
   assign  s_logisimBus47[32]  =  1'b0;
   assign  s_logisimBus47[33]  =  1'b0;
   assign  s_logisimBus47[34]  =  1'b0;
   assign  s_logisimBus47[35]  =  1'b0;
   assign  s_logisimBus47[36]  =  1'b0;
   assign  s_logisimBus47[37]  =  1'b0;
   assign  s_logisimBus47[38]  =  1'b0;
   assign  s_logisimBus47[39]  =  1'b0;
   assign  s_logisimBus47[40]  =  1'b0;
   assign  s_logisimBus47[41]  =  1'b0;
   assign  s_logisimBus47[42]  =  1'b0;
   assign  s_logisimBus47[43]  =  1'b0;
   assign  s_logisimBus47[44]  =  1'b0;
   assign  s_logisimBus47[45]  =  1'b0;
   assign  s_logisimBus47[46]  =  1'b0;
   assign  s_logisimBus47[47]  =  1'b0;
   assign  s_logisimBus47[48]  =  1'b0;
   assign  s_logisimBus47[49]  =  1'b0;
   assign  s_logisimBus47[50]  =  1'b0;
   assign  s_logisimBus47[51]  =  1'b0;
   assign  s_logisimBus47[52]  =  1'b0;
   assign  s_logisimBus47[53]  =  1'b0;
   assign  s_logisimBus47[54]  =  1'b0;
   assign  s_logisimBus47[55]  =  1'b0;
   assign  s_logisimBus47[56]  =  1'b0;
   assign  s_logisimBus47[57]  =  1'b0;
   assign  s_logisimBus47[58]  =  1'b0;
   assign  s_logisimBus47[59]  =  1'b0;
   assign  s_logisimBus47[60]  =  1'b0;
   assign  s_logisimBus47[61]  =  1'b0;
   assign  s_logisimBus47[62]  =  1'b0;
   assign  s_logisimBus47[63]  =  1'b0;


   // Constant
   assign  s_logisimBus23[30:0]  =  {3'b111, 28'hF800000};


   // Constant
   assign  s_logisimBus119[7:0]  =  8'h01;


   // Constant
   assign  s_logisimBus80[30:0]  =  {3'b111, 28'hFC00000};


   // NOT Gate
   assign s_logisimNet145 = ~s_logisimNet51;

   // NOT Gate
   assign s_logisimNet55 = ~s_logisimNet95;

   // NOT Gate
   assign s_logisimNet30 = ~s_logisimNet152;

   /*******************************************************************************
   ** Here all normal components are defined                                     **
   *******************************************************************************/
   AND_GATE #(.BubblesMask(2'b00))
      GATES_1 (.input1(s_logisimNet15),
               .input2(s_logisimNet130),
               .result(s_logisimNet2));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_2 (.input1(s_logisimNet74),
               .input2(s_logisimNet125),
               .result(s_logisimNet45));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_3 (.input1(s_logisimNet0),
               .input2(s_logisimNet79),
               .result(s_logisimNet96));

   OR_GATE_3_INPUTS #(.BubblesMask(3'b000))
      GATES_4 (.input1(s_logisimNet96),
               .input2(s_logisimNet45),
               .input3(s_logisimNet2),
               .result(s_logisimNet10));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_5 (.input1(s_logisimNet121),
               .input2(s_logisimNet159),
               .result(s_logisimNet8));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_6 (.input1(s_logisimNet70),
               .input2(s_logisimNet158),
               .result(s_logisimNet122));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_7 (.input1(s_logisimNet102),
               .input2(s_logisimNet145),
               .result(s_logisimNet81));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_8 (.input1(s_logisimNet64),
               .input2(s_logisimNet76),
               .result(s_logisimNet44));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_9 (.input1(s_logisimNet38),
               .input2(s_logisimNet55),
               .result(s_logisimNet19));

   AND_GATE #(.BubblesMask(2'b00))
      GATES_10 (.input1(s_logisimNet62),
                .input2(s_logisimNet112),
                .result(s_logisimNet66));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_11 (.input1(s_logisimNet19),
                .input2(s_logisimNet81),
                .result(s_logisimNet129));

   OR_GATE #(.BubblesMask(2'b00))
      GATES_12 (.input1(s_logisimNet66),
                .input2(s_logisimNet44),
                .result(s_logisimNet105));

   Multiplexer_bus_2 #(.nrOfBits(32))
      PLEXERS_13 (.enable(1'b1),
                  .muxIn_0(s_logisimBus94[31:0]),
                  .muxIn_1(s_logisimBus23[31:0]),
                  .muxOut(s_logisimBus115[31:0]),
                  .sel(s_logisimNet105));

   Multiplexer_bus_2 #(.nrOfBits(32))
      PLEXERS_14 (.enable(1'b1),
                  .muxIn_0(s_logisimBus115[31:0]),
                  .muxIn_1(s_logisimBus80[31:0]),
                  .muxOut(s_logisimBus24[31:0]),
                  .sel(s_logisimNet129));

   Multiplexer_2   PLEXERS_15 (.enable(1'b1),
                               .muxIn_0(s_logisimNet124),
                               .muxIn_1(s_logisimBus43[1]),
                               .muxOut(s_logisimNet130),
                               .sel(s_logisimBus27[23]));

   Multiplexer_bus_2 #(.nrOfBits(8))
      PLEXERS_16 (.enable(1'b1),
                  .muxIn_0(s_logisimBus36[7:0]),
                  .muxIn_1(s_logisimBus6[7:0]),
                  .muxOut(s_logisimBus32[30:23]),
                  .sel(s_logisimNet10));

   Multiplexer_bus_2 #(.nrOfBits(23))
      PLEXERS_17 (.enable(1'b1),
                  .muxIn_0(s_logisimBus149[22:0]),
                  .muxIn_1(s_logisimBus20[22:0]),
                  .muxOut(s_logisimBus68[22:0]),
                  .sel(s_logisimNet130));

   Multiplexer_2   PLEXERS_18 (.enable(1'b1),
                               .muxIn_0(s_logisimNet118),
                               .muxIn_1(s_logisimNet56),
                               .muxOut(s_logisimNet121),
                               .sel(s_logisimNet21));

   Multiplexer_2   PLEXERS_19 (.enable(1'b1),
                               .muxIn_0(s_logisimNet46),
                               .muxIn_1(s_logisimNet7),
                               .muxOut(s_logisimNet70),
                               .sel(s_logisimNet92));

   Multiplexer_bus_2 #(.nrOfBits(23))
      PLEXERS_20 (.enable(1'b1),
                  .muxIn_0(s_logisimBus108[22:0]),
                  .muxIn_1(s_logisimBus34[22:0]),
                  .muxOut(s_logisimBus83[22:0]),
                  .sel(s_logisimNet79));

   Multiplexer_bus_2 #(.nrOfBits(23))
      PLEXERS_21 (.enable(1'b1),
                  .muxIn_0(s_logisimBus142[22:0]),
                  .muxIn_1(s_logisimBus58[22:0]),
                  .muxOut(s_logisimBus50[22:0]),
                  .sel(s_logisimNet125));

   Multiplexer_bus_2 #(.nrOfBits(23))
      PLEXERS_22 (.enable(1'b1),
                  .muxIn_0(s_logisimBus83[22:0]),
                  .muxIn_1(s_logisimBus3[22:0]),
                  .muxOut(s_logisimBus126[22:0]),
                  .sel(s_logisimNet8));

   Multiplexer_bus_2 #(.nrOfBits(23))
      PLEXERS_23 (.enable(1'b1),
                  .muxIn_0(s_logisimBus50[22:0]),
                  .muxIn_1(s_logisimBus117[22:0]),
                  .muxOut(s_logisimBus100[22:0]),
                  .sel(s_logisimNet122));

   Multiplexer_bus_2 #(.nrOfBits(32))
      PLEXERS_24 (.enable(1'b1),
                  .muxIn_0(s_logisimBus61[31:0]),
                  .muxIn_1(s_logisimBus53[31:0]),
                  .muxOut(s_logisimBus103[31:0]),
                  .sel(s_logisimBus4[23]));

   Multiplexer_bus_2 #(.nrOfBits(32))
      PLEXERS_25 (.enable(1'b1),
                  .muxIn_0(s_logisimBus106[31:0]),
                  .muxIn_1(s_logisimBus1[31:0]),
                  .muxOut(s_logisimBus89[31:0]),
                  .sel(s_logisimBus27[23]));

   Multiplexer_2   PLEXERS_26 (.enable(1'b1),
                               .muxIn_0(s_logisimNet116),
                               .muxIn_1(s_logisimNet67),
                               .muxOut(s_logisimBus27[23]),
                               .sel(s_logisimNet17));

   Multiplexer_2   PLEXERS_27 (.enable(1'b1),
                               .muxIn_0(s_logisimNet59),
                               .muxIn_1(s_logisimNet139),
                               .muxOut(s_logisimBus4[23]),
                               .sel(s_logisimNet26));

   Multiplexer_2   PLEXERS_28 (.enable(1'b1),
                               .muxIn_0(s_logisimBus134[31]),
                               .muxIn_1(s_logisimNet156),
                               .muxOut(s_logisimBus23[31]),
                               .sel(s_logisimNet66));

   Multiplexer_2   PLEXERS_29 (.enable(1'b1),
                               .muxIn_0(s_logisimBus134[31]),
                               .muxIn_1(s_logisimNet156),
                               .muxOut(s_logisimBus80[31]),
                               .sel(s_logisimNet19));

   Multiplexer_bus_2 #(.nrOfBits(32))
      PLEXERS_30 (.enable(1'b1),
                  .muxIn_0(s_logisimBus32[31:0]),
                  .muxIn_1(s_logisimBus133[31:0]),
                  .muxOut(s_logisimBus94[31:0]),
                  .sel(s_logisimNet30));

   Multiplexer_bus_2 #(.nrOfBits(23))
      PLEXERS_31 (.enable(1'b1),
                  .muxIn_0(s_logisimBus126[22:0]),
                  .muxIn_1(s_logisimBus100[22:0]),
                  .muxOut(s_logisimBus147[22:0]),
                  .sel(s_logisimNet73));

   Multiplexer_bus_2 #(.nrOfBits(8))
      PLEXERS_32 (.enable(1'b1),
                  .muxIn_0(s_logisimBus140[7:0]),
                  .muxIn_1(s_logisimBus151[7:0]),
                  .muxOut(s_logisimBus36[7:0]),
                  .sel(s_logisimNet0));

   Multiplexer_bus_2 #(.nrOfBits(23))
      PLEXERS_33 (.enable(1'b1),
                  .muxIn_0(s_logisimBus149[22:0]),
                  .muxIn_1(s_logisimBus101[22:0]),
                  .muxOut(s_logisimBus20[22:0]),
                  .sel(s_logisimBus27[23]));

   Multiplexer_bus_2 #(.nrOfBits(23))
      PLEXERS_34 (.enable(1'b1),
                  .muxIn_0(s_logisimBus147[22:0]),
                  .muxIn_1(s_logisimBus68[22:0]),
                  .muxOut(s_logisimBus32[22:0]),
                  .sel(s_logisimNet16));

   Comparator #(.nrOfBits(32),
                .twosComplement(1))
      ARITH_35 (.aEqualsB(),
                .aGreaterThanB(),
                .aLessThanB(s_logisimNet21),
                .dataA(s_logisimBus103[31:0]),
                .dataB(s_logisimBus146[31:0]));

   Shifter_23_bit #(.shifterMode(2))
      ARITH_36 (.dataA(s_logisimBus108[22:0]),
                .result(s_logisimBus34[22:0]),
                .shiftAmount(s_logisimBus91[4:0]));

   Shifter_23_bit #(.shifterMode(2))
      ARITH_37 (.dataA(s_logisimBus142[22:0]),
                .result(s_logisimBus58[22:0]),
                .shiftAmount(s_logisimBus33[4:0]));

   Subtractor #(.extendedBits(10),
                .nrOfBits(9))
      ARITH_38 (.borrowIn(1'b0),
                .borrowOut(),
                .dataA(s_logisimBus35[8:0]),
                .dataB(s_logisimBus22[8:0]),
                .result(s_logisimBus60[8:0]));

   Subtractor #(.extendedBits(10),
                .nrOfBits(9))
      ARITH_39 (.borrowIn(1'b0),
                .borrowOut(),
                .dataA(s_logisimBus48[8:0]),
                .dataB(s_logisimBus69[8:0]),
                .result(s_logisimBus14[8:0]));

   Comparator #(.nrOfBits(32),
                .twosComplement(1))
      ARITH_40 (.aEqualsB(),
                .aGreaterThanB(),
                .aLessThanB(s_logisimNet92),
                .dataA(s_logisimBus89[31:0]),
                .dataB(s_logisimBus75[31:0]));

   Comparator #(.nrOfBits(9),
                .twosComplement(1))
      ARITH_41 (.aEqualsB(),
                .aGreaterThanB(),
                .aLessThanB(),
                .dataA(s_logisimBus60[8:0]),
                .dataB(s_logisimBus131[8:0]));

   Comparator #(.nrOfBits(9),
                .twosComplement(1))
      ARITH_42 (.aEqualsB(),
                .aGreaterThanB(),
                .aLessThanB(),
                .dataA(s_logisimBus14[8:0]),
                .dataB(s_logisimBus107[8:0]));

   Adder #(.extendedBits(24),
           .nrOfBits(23))
      ARITH_43 (.carryIn(1'b0),
                .carryOut(),
                .dataA(s_logisimBus83[22:0]),
                .dataB(s_logisimBus128[22:0]),
                .result(s_logisimBus3[22:0]));

   Subtractor #(.extendedBits(9),
                .nrOfBits(8))
      ARITH_44 (.borrowIn(1'b0),
                .borrowOut(),
                .dataA(s_logisimBus140[7:0]),
                .dataB(s_logisimBus151[7:0]),
                .result(s_logisimBus137[7:0]));

   Adder #(.extendedBits(24),
           .nrOfBits(23))
      ARITH_45 (.carryIn(1'b0),
                .carryOut(),
                .dataA(s_logisimBus50[22:0]),
                .dataB(s_logisimBus104[22:0]),
                .result(s_logisimBus117[22:0]));

   Subtractor #(.extendedBits(9),
                .nrOfBits(8))
      ARITH_46 (.borrowIn(1'b0),
                .borrowOut(),
                .dataA(s_logisimBus151[7:0]),
                .dataB(s_logisimBus140[7:0]),
                .result(s_logisimBus97[7:0]));

   Subtractor #(.extendedBits(33),
                .nrOfBits(32))
      ARITH_47 (.borrowIn(1'b0),
                .borrowOut(),
                .dataA(s_logisimBus53[31:0]),
                .dataB(s_logisimBus110[31:0]),
                .result(s_logisimBus61[31:0]));

   Subtractor #(.extendedBits(33),
                .nrOfBits(32))
      ARITH_48 (.borrowIn(1'b0),
                .borrowOut(),
                .dataA(s_logisimBus1[31:0]),
                .dataB(s_logisimBus153[31:0]),
                .result(s_logisimBus106[31:0]));

   Adder #(.extendedBits(24),
           .nrOfBits(23))
      ARITH_49 (.carryIn(1'b0),
                .carryOut(s_logisimNet124),
                .dataA(s_logisimBus148[22:0]),
                .dataB(s_logisimBus135[22:0]),
                .result(s_logisimBus149[22:0]));

   Comparator #(.nrOfBits(23),
                .twosComplement(1))
      ARITH_50 (.aEqualsB(s_logisimNet51),
                .aGreaterThanB(),
                .aLessThanB(),
                .dataA(s_logisimBus148[22:0]),
                .dataB(s_logisimBus114[22:0]));

   Comparator #(.nrOfBits(23),
                .twosComplement(1))
      ARITH_51 (.aEqualsB(s_logisimNet76),
                .aGreaterThanB(),
                .aLessThanB(),
                .dataA(s_logisimBus148[22:0]),
                .dataB(s_logisimBus85[22:0]));

   Comparator #(.nrOfBits(23),
                .twosComplement(1))
      ARITH_52 (.aEqualsB(s_logisimNet95),
                .aGreaterThanB(),
                .aLessThanB(),
                .dataA(s_logisimBus135[22:0]),
                .dataB(s_logisimBus12[22:0]));

   Comparator #(.nrOfBits(8),
                .twosComplement(1))
      ARITH_53 (.aEqualsB(s_logisimNet102),
                .aGreaterThanB(),
                .aLessThanB(),
                .dataA(s_logisimBus140[7:0]),
                .dataB(s_logisimBus37[7:0]));

   Comparator #(.nrOfBits(23),
                .twosComplement(1))
      ARITH_54 (.aEqualsB(s_logisimNet112),
                .aGreaterThanB(),
                .aLessThanB(),
                .dataA(s_logisimBus135[22:0]),
                .dataB(s_logisimBus123[22:0]));

   Comparator #(.nrOfBits(8),
                .twosComplement(1))
      ARITH_55 (.aEqualsB(s_logisimNet64),
                .aGreaterThanB(),
                .aLessThanB(),
                .dataA(s_logisimBus140[7:0]),
                .dataB(s_logisimBus136[7:0]));

   Comparator #(.nrOfBits(8),
                .twosComplement(1))
      ARITH_56 (.aEqualsB(s_logisimNet38),
                .aGreaterThanB(),
                .aLessThanB(),
                .dataA(s_logisimBus151[7:0]),
                .dataB(s_logisimBus84[7:0]));

   Comparator #(.nrOfBits(8),
                .twosComplement(1))
      ARITH_57 (.aEqualsB(s_logisimNet62),
                .aGreaterThanB(),
                .aLessThanB(),
                .dataA(s_logisimBus151[7:0]),
                .dataB(s_logisimBus49[7:0]));

   Adder #(.extendedBits(3),
           .nrOfBits(2))
      ARITH_58 (.carryIn(1'b0),
                .carryOut(),
                .dataA(s_logisimBus13[1:0]),
                .dataB(s_logisimBus109[1:0]),
                .result(s_logisimBus43[1:0]));

   Comparator #(.nrOfBits(8),
                .twosComplement(1))
      ARITH_59 (.aEqualsB(s_logisimNet17),
                .aGreaterThanB(),
                .aLessThanB(),
                .dataA(s_logisimBus140[7:0]),
                .dataB(s_logisimBus150[7:0]));

   Comparator #(.nrOfBits(8),
                .twosComplement(1))
      ARITH_60 (.aEqualsB(s_logisimNet26),
                .aGreaterThanB(),
                .aLessThanB(),
                .dataA(s_logisimBus151[7:0]),
                .dataB(s_logisimBus93[7:0]));

   BitComparator #(.twosComplement(1))
      ARITH_61 (.aEqualsB(s_logisimNet152),
                .aGreaterThanB(),
                .aLessThanB(),
                .dataA(s_logisimNet156),
                .dataB(s_logisimBus134[31]));

   Comparator #(.nrOfBits(9),
                .twosComplement(1))
      ARITH_62 (.aEqualsB(s_logisimNet16),
                .aGreaterThanB(s_logisimNet73),
                .aLessThanB(),
                .dataA(s_logisimBus5[8:0]),
                .dataB(s_logisimBus87[8:0]));

   Subtractor #(.extendedBits(33),
                .nrOfBits(32))
      ARITH_63 (.borrowIn(1'b0),
                .borrowOut(),
                .dataA(s_logisimBus9[31:0]),
                .dataB(s_logisimBus144[31:0]),
                .result(s_logisimBus52[31:0]));

   Comparator #(.nrOfBits(9),
                .twosComplement(1))
      ARITH_64 (.aEqualsB(s_logisimNet15),
                .aGreaterThanB(s_logisimNet0),
                .aLessThanB(s_logisimNet74),
                .dataA(s_logisimBus88[8:0]),
                .dataB(s_logisimBus29[8:0]));

   Subtractor #(.extendedBits(33),
                .nrOfBits(32))
      ARITH_65 (.borrowIn(1'b0),
                .borrowOut(),
                .dataA(s_logisimBus11[31:0]),
                .dataB(s_logisimBus132[31:0]),
                .result(s_logisimBus57[31:0]));

   Adder #(.extendedBits(24),
           .nrOfBits(23))
      ARITH_66 (.carryIn(1'b0),
                .carryOut(s_logisimNet25),
                .dataA(s_logisimBus42[22:0]),
                .dataB(s_logisimBus148[22:0]),
                .result(s_logisimBus108[22:0]));

   Adder #(.extendedBits(24),
           .nrOfBits(23))
      ARITH_67 (.carryIn(1'b0),
                .carryOut(s_logisimNet65),
                .dataA(s_logisimBus78[22:0]),
                .dataB(s_logisimBus135[22:0]),
                .result(s_logisimBus142[22:0]));

   FullAdder #(.extendedBits(2))
      ARITH_68 (.carryIn(1'b0),
                .carryOut(s_logisimNet79),
                .dataA(s_logisimNet25),
                .dataB(s_logisimBus27[23]),
                .result());

   FullAdder #(.extendedBits(2))
      ARITH_69 (.carryIn(1'b0),
                .carryOut(s_logisimNet125),
                .dataA(s_logisimNet65),
                .dataB(s_logisimBus4[23]),
                .result());

   Adder #(.extendedBits(9),
           .nrOfBits(8))
      ARITH_70 (.carryIn(1'b0),
                .carryOut(),
                .dataA(s_logisimBus36[7:0]),
                .dataB(s_logisimBus119[7:0]),
                .result(s_logisimBus6[7:0]));


   /*******************************************************************************
   ** Here all sub-circuits are defined                                          **
   *******************************************************************************/

   add_find_bit_1   v29 (.number(s_logisimBus47[63:0]),
                         .s(s_logisimNet7),
                         .shift(s_logisimBus89[5:0]),
                         .sticky(s_logisimNet158));

   fMinnus   v23 (.a(s_logisimBus127[31:0]),
                  .b(s_logisimBus134[31:0]),
                  .res(s_logisimBus133[31:0]));

   SRL_fadd   v24 (.a(s_logisimBus9[31:0]),
                   .b(s_logisimBus103[31:0]),
                   .one_signal(),
                   .res_low(s_logisimBus42[31:0]));

   SRL_fadd   v27 (.a(s_logisimBus11[31:0]),
                   .b(s_logisimBus89[31:0]),
                   .one_signal(),
                   .res_low(s_logisimBus78[31:0]));

   SLLL   v25 (.a(s_logisimBus42[31:0]),
               .b(s_logisimBus103[31:0]),
               .res_high(),
               .res_low(s_logisimBus144[31:0]));

   SLLL   v28 (.a(s_logisimBus78[31:0]),
               .b(s_logisimBus89[31:0]),
               .res_high(),
               .res_low(s_logisimBus132[31:0]));

   add_find_bit_1   v26 (.number(s_logisimBus82[63:0]),
                         .s(s_logisimNet56),
                         .shift(s_logisimBus103[5:0]),
                         .sticky(s_logisimNet159));

endmodule
