/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
CU5
**
**
**
*****************************************************************************/
module
CU5(
func,
link,
memToReg,
opCode,
regWrite
);
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
[5:0]
func;
input
[5:0]
opCode;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
link;
output
memToReg;
output
regWrite;
/*******************************************************************************
**
The
wires
are
defined
here
**
*******************************************************************************/
wire
[3:0]
s_logisimBus10;
wire
[3:0]
s_logisimBus11;
wire
[3:0]
s_logisimBus12;
wire
[3:0]
s_logisimBus13;
wire
[3:0]
s_logisimBus20;
wire
[3:0]
s_logisimBus21;
wire
[3:0]
s_logisimBus24;
wire
[3:0]
s_logisimBus26;
wire
[3:0]
s_logisimBus27;
wire
[3:0]
s_logisimBus39;
wire
[3:0]
s_logisimBus40;
wire
[3:0]
s_logisimBus41;
wire
[3:0]
s_logisimBus42;
wire
[3:0]
s_logisimBus43;
wire
[3:0]
s_logisimBus44;
wire
[3:0]
s_logisimBus45;
wire
[3:0]
s_logisimBus46;
wire
[3:0]
s_logisimBus47;
wire
[3:0]
s_logisimBus48;
wire
[3:0]
s_logisimBus49;
wire
[5:0]
s_logisimBus5;
wire
[3:0]
s_logisimBus50;
wire
[3:0]
s_logisimBus51;
wire
[5:0]
s_logisimBus52;
wire
[5:0]
s_logisimBus54;
wire
[5:0]
s_logisimBus55;
wire
[5:0]
s_logisimBus56;
wire
[5:0]
s_logisimBus57;
wire
[5:0]
s_logisimBus58;
wire
[5:0]
s_logisimBus59;
wire
[5:0]
s_logisimBus6;
wire
[5:0]
s_logisimBus60;
wire
[5:0]
s_logisimBus61;
wire
[5:0]
s_logisimBus62;
wire
[5:0]
s_logisimBus63;
wire
[5:0]
s_logisimBus64;
wire
[5:0]
s_logisimBus65;
wire
[5:0]
s_logisimBus66;
wire
[5:0]
s_logisimBus67;
wire
[5:0]
s_logisimBus68;
wire
[5:0]
s_logisimBus69;
wire
[3:0]
s_logisimBus7;
wire
[5:0]
s_logisimBus70;
wire
[5:0]
s_logisimBus71;
wire
[5:0]
s_logisimBus72;
wire
[5:0]
s_logisimBus73;
wire
[5:0]
s_logisimBus74;
wire
[5:0]
s_logisimBus75;
wire
[5:0]
s_logisimBus76;
wire
[3:0]
s_logisimBus8;
wire
s_logisimNet0;
wire
s_logisimNet1;
wire
s_logisimNet14;
wire
s_logisimNet15;
wire
s_logisimNet16;
wire
s_logisimNet17;
wire
s_logisimNet18;
wire
s_logisimNet19;
wire
s_logisimNet2;
wire
s_logisimNet22;
wire
s_logisimNet23;
wire
s_logisimNet25;
wire
s_logisimNet28;
wire
s_logisimNet29;
wire
s_logisimNet3;
wire
s_logisimNet30;
wire
s_logisimNet31;
wire
s_logisimNet32;
wire
s_logisimNet33;
wire
s_logisimNet34;
wire
s_logisimNet35;
wire
s_logisimNet36;
wire
s_logisimNet37;
wire
s_logisimNet38;
wire
s_logisimNet4;
wire
s_logisimNet53;
wire
s_logisimNet9;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
/*******************************************************************************
**
Here
all
input
connections
are
defined
**
*******************************************************************************/
assign
s_logisimBus5[5:0]
=
opCode;
assign
s_logisimBus6[5:0]
=
func;
/*******************************************************************************
**
Here
all
output
connections
are
defined
**
*******************************************************************************/
assign
link
=
s_logisimNet18;
assign
memToReg
=
s_logisimNet35;
assign
regWrite
=
s_logisimNet28;
/*******************************************************************************
**
Here
all
in-lined
components
are
defined
**
*******************************************************************************/
assign
s_logisimBus52[5:0]
=
{2'b10,
4'h0};
assign
s_logisimBus54[5:0]
=
{2'b10,
4'h2};
assign
s_logisimBus55[5:0]
=
{2'b10,
4'h4};
assign
s_logisimBus56[5:0]
=
{2'b10,
4'h5};
assign
s_logisimBus57[5:0]
=
{2'b10,
4'h6};
assign
s_logisimBus58[5:0]
=
{2'b00,
4'h4};
assign
s_logisimBus59[5:0]
=
{2'b00,
4'h6};
assign
s_logisimBus60[5:0]
=
{2'b00,
4'h7};
assign
s_logisimBus61[5:0]
=
{2'b01,
4'hA};
assign
s_logisimBus62[5:0]
=
{2'b01,
4'h0};
assign
s_logisimBus63[5:0]
=
{2'b00,
4'h0};
assign
s_logisimBus64[5:0]
=
{2'b00,
4'h8};
assign
s_logisimBus65[5:0]
=
{2'b01,
4'h2};
assign
s_logisimBus66[5:0]
=
{2'b00,
4'h2};
assign
s_logisimBus39[3:0]
=
4'h0;
assign
s_logisimBus40[3:0]
=
4'h1;
assign
s_logisimBus41[3:0]
=
4'h4;
assign
s_logisimBus42[3:0]
=
4'h5;
assign
s_logisimBus43[3:0]
=
4'h6;
assign
s_logisimBus67[5:0]
=
{2'b00,
4'h0};
assign
s_logisimBus68[5:0]
=
{2'b00,
4'h8};
assign
s_logisimBus69[5:0]
=
{2'b10,
4'hB};
assign
s_logisimBus70[5:0]
=
{2'b10,
4'h3};
assign
s_logisimBus71[5:0]
=
{2'b00,
4'h5};
assign
s_logisimBus72[5:0]
=
{2'b00,
4'hA};
assign
s_logisimBus73[5:0]
=
{2'b00,
4'h2};
assign
s_logisimBus74[5:0]
=
{2'b00,
4'h3};
assign
s_logisimBus75[5:0]
=
{2'b00,
4'h4};
assign
s_logisimBus76[5:0]
=
{2'b01,
4'hC};
assign
s_logisimBus44[3:0]
=
4'h9;
assign
s_logisimBus45[3:0]
=
4'hA;
assign
s_logisimBus46[3:0]
=
4'hB;
assign
s_logisimBus47[3:0]
=
4'h3;
assign
s_logisimBus48[3:0]
=
4'hF;
assign
s_logisimBus49[3:0]
=
4'h9;
assign
s_logisimBus50[3:0]
=
4'hF;
assign
s_logisimBus51[3:0]
=
4'hF;
/*******************************************************************************
**
Here
all
normal
components
are
defined
**
*******************************************************************************/
AND_GATE
#(.BubblesMask(2'b01))
GATES_1
(.input1(s_logisimNet17),
.input2(s_logisimNet31),
.result(s_logisimNet3));
AND_GATE
#(.BubblesMask(2'b00))
GATES_2
(.input1(s_logisimNet2),
.input2(s_logisimNet38),
.result(s_logisimNet37));
OR_GATE_5_INPUTS
#(.BubblesMask({1'b0,
4'h0}))
GATES_3
(.input1(s_logisimNet3),
.input2(s_logisimNet25),
.input3(s_logisimNet37),
.input4(s_logisimNet36),
.input5(s_logisimNet35),
.result(s_logisimNet28));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_4
(.enable(1'b1),
.muxIn_0(s_logisimBus39[3:0]),
.muxIn_1(s_logisimBus40[3:0]),
.muxOut(s_logisimBus8[3:0]),
.sel(s_logisimNet19));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_5
(.enable(1'b1),
.muxIn_0(s_logisimBus8[3:0]),
.muxIn_1(s_logisimBus41[3:0]),
.muxOut(s_logisimBus7[3:0]),
.sel(s_logisimNet15));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_6
(.enable(1'b1),
.muxIn_0(s_logisimBus7[3:0]),
.muxIn_1(s_logisimBus42[3:0]),
.muxOut(s_logisimBus27[3:0]),
.sel(s_logisimNet0));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_7
(.enable(1'b1),
.muxIn_0(s_logisimBus27[3:0]),
.muxIn_1(s_logisimBus43[3:0]),
.muxOut(s_logisimBus21[3:0]),
.sel(s_logisimNet29));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_8
(.enable(1'b1),
.muxIn_0(s_logisimBus21[3:0]),
.muxIn_1(s_logisimBus44[3:0]),
.muxOut(s_logisimBus11[3:0]),
.sel(s_logisimNet23));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_9
(.enable(1'b1),
.muxIn_0(s_logisimBus11[3:0]),
.muxIn_1(s_logisimBus45[3:0]),
.muxOut(s_logisimBus13[3:0]),
.sel(s_logisimNet4));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_10
(.enable(1'b1),
.muxIn_0(s_logisimBus13[3:0]),
.muxIn_1(s_logisimBus46[3:0]),
.muxOut(s_logisimBus26[3:0]),
.sel(s_logisimNet1));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_11
(.enable(1'b1),
.muxIn_0(s_logisimBus26[3:0]),
.muxIn_1(s_logisimBus47[3:0]),
.muxOut(s_logisimBus20[3:0]),
.sel(s_logisimNet16));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_12
(.enable(1'b1),
.muxIn_0(s_logisimBus20[3:0]),
.muxIn_1(s_logisimBus48[3:0]),
.muxOut(s_logisimBus10[3:0]),
.sel(s_logisimNet22));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_13
(.enable(1'b1),
.muxIn_0(s_logisimBus10[3:0]),
.muxIn_1(s_logisimBus49[3:0]),
.muxOut(s_logisimBus12[3:0]),
.sel(s_logisimNet14));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_14
(.enable(1'b1),
.muxIn_0(s_logisimBus12[3:0]),
.muxIn_1(s_logisimBus50[3:0]),
.muxOut(s_logisimBus24[3:0]),
.sel(s_logisimNet17));
Multiplexer_bus_2
#(.nrOfBits(4))
PLEXERS_15
(.enable(1'b1),
.muxIn_0(s_logisimBus24[3:0]),
.muxIn_1(s_logisimBus51[3:0]),
.muxOut(),
.sel(s_logisimNet9));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_16
(.aEqualsB(s_logisimNet53),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus52[5:0]),
.dataB(s_logisimBus6[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_17
(.aEqualsB(s_logisimNet19),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus54[5:0]),
.dataB(s_logisimBus6[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_18
(.aEqualsB(s_logisimNet15),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus55[5:0]),
.dataB(s_logisimBus6[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_19
(.aEqualsB(s_logisimNet0),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus56[5:0]),
.dataB(s_logisimBus6[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_20
(.aEqualsB(s_logisimNet29),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus57[5:0]),
.dataB(s_logisimBus6[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_21
(.aEqualsB(s_logisimNet23),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus58[5:0]),
.dataB(s_logisimBus6[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_22
(.aEqualsB(s_logisimNet4),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus59[5:0]),
.dataB(s_logisimBus6[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_23
(.aEqualsB(s_logisimNet1),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus60[5:0]),
.dataB(s_logisimBus6[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_24
(.aEqualsB(s_logisimNet16),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus61[5:0]),
.dataB(s_logisimBus6[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_25
(.aEqualsB(s_logisimNet22),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus62[5:0]),
.dataB(s_logisimBus6[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_26
(.aEqualsB(s_logisimNet14),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus63[5:0]),
.dataB(s_logisimBus6[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_27
(.aEqualsB(s_logisimNet17),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus64[5:0]),
.dataB(s_logisimBus6[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_28
(.aEqualsB(s_logisimNet9),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus65[5:0]),
.dataB(s_logisimBus6[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_29
(.aEqualsB(s_logisimNet38),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus66[5:0]),
.dataB(s_logisimBus6[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_30
(.aEqualsB(s_logisimNet31),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus67[5:0]),
.dataB(s_logisimBus5[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_31
(.aEqualsB(s_logisimNet25),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus68[5:0]),
.dataB(s_logisimBus5[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_32
(.aEqualsB(s_logisimNet30),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus69[5:0]),
.dataB(s_logisimBus5[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_33
(.aEqualsB(s_logisimNet35),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus70[5:0]),
.dataB(s_logisimBus5[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_34
(.aEqualsB(s_logisimNet32),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus71[5:0]),
.dataB(s_logisimBus5[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_35
(.aEqualsB(s_logisimNet36),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus72[5:0]),
.dataB(s_logisimBus5[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_36
(.aEqualsB(s_logisimNet33),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus73[5:0]),
.dataB(s_logisimBus5[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_37
(.aEqualsB(s_logisimNet18),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus74[5:0]),
.dataB(s_logisimBus5[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_38
(.aEqualsB(s_logisimNet34),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus75[5:0]),
.dataB(s_logisimBus5[5:0]));
Comparator
#(.nrOfBits(6),
.twosComplement(0))
ARITH_39
(.aEqualsB(s_logisimNet2),
.aGreaterThanB(),
.aLessThanB(),
.dataA(s_logisimBus76[5:0]),
.dataB(s_logisimBus5[5:0]));
endmodule