/******************************************************************************
**
Logisim-evolution
goes
FPGA
automatic
generated
Verilog
code
**
**
https://github.com/logisim-evolution/
**
**
**
**
Component
:
Negator
**
**
**
*****************************************************************************/
module
Negator(
dataX,
minDataX
);
/*******************************************************************************
**
Here
all
module
parameters
are
defined
with
a
dummy
value
**
*******************************************************************************/
parameter
nrOfBits
=
1;
/*******************************************************************************
**
The
inputs
are
defined
here
**
*******************************************************************************/
input
[nrOfBits-1:0]
dataX;
/*******************************************************************************
**
The
outputs
are
defined
here
**
*******************************************************************************/
output
[nrOfBits-1:0]
minDataX;
/*******************************************************************************
**
The
module
functionality
is
described
here
**
*******************************************************************************/
assign
minDataX
=
-dataX;
endmodule